��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�UΣ<iZB\���@s�Pg�eW��t!����߬ �j,�k�
B���R/�;��	���{���Gx�e���
+�-�)2�q����8�Z�E�3`p��,�Vh5"�]6���Qm@I�1��ܟ��UU�	�$��5��~������ܠ����LG���X1���A<` v5�
���a��K�ZT����һ�����̀3�\�p1.�OJ���Bªu���dW�f�]O��^�/�*PɞI�o�l�C��93Nʼy��a��E"t�e��ށ��;@,��FH�A� �\�\�1/���_���?��/� Qk0^�ƥ�iO�Z�O�Ϸ���~R�5h���	��4��ٺQ�Ϭ�|a&�� ���0ÌM�L�fV����%�*3�В���������#���ɱ�m� 7��/z���/v�4�6GTN�p�^v���-p�y�*С�ϳDyl;03�<cG�����6T��(2�J!�&������o��pa��I���n��މ�����W3�F�BB��aR�J� koq���h�rTH��7�JZ�L)ݽ�|u ��u�
��E��g6�G/�,:v��iS�Ƙl��:�r=7� ��]�w�=2l�G2h`騤��C�K��zCA�S^�B�sC�;�
O�d䟪=�v7-�����?<� ��[��6A�k9���q�Mx�4y�/2�01������l�Tx�������s�@���
�.�e"���()�@,�,+��m��!��*w�� A�q|D���Qd��#���!�L�$-�ǌ��L)X�.�������r���>� ,�ɂ����pӄ�U�Mx6]���E!�敢p���}&�\08"Xgg��fN���*� ����J/���	�$;#@U殶]A�E�XI��vﵒ�B�i�	�8��"/�}s�:8_>�܈+m}8t 1P�P�؟hyQ5�ʳU��v����e���(�*��W�����b}�0���	��]��0L�4!'@�S��L,�;����@.�{�j�����[i�O��Y���^�}�ƻׁ\��<z�@���[{��_�% ���n�٤`�)���U�����G�V����Y�Ϊ�zrJmN���r�Xe~q�*�y�}Gi7�𑢵LMl|�,����d��*&�!D��T�l厄? I�"h�i�ߺ�`�7�(�:`1�L�t�H���D,���x���*�q�Q�zc��_[<X�NR�	kʑ?��we%�����<oߛ��/�H݁K�lJ5 FyM���Ԍ-�9�c�[�2�t��A2U��2*)SތS�&�&Ӎ���K\�Q��;_:�~f����N5��U�~�p2Q��'�3��h�W�TslK�N ]�xig�hp��p�Uk3��k@P��>����
"1��4��ëQ3K��f��*+ae���Z�`�vQ�C9�
��d'`N��d5��g5���=��'l �oB� W."G�A�E�D�ál��A�tW=<T{1p���T.Ţ4�@��[��O����r܎���D,��������ܙ�c�@=׋�S�\�
7ԟ��yS��̧W��~	 ��L�L��@���0mƿr�tb1@���N������B<�� 3n�I�]�w�R@+3݇�����~{����(��j.�,E���O���Nf�4"�u��J��jڍt;�Q�Þ��+C \5�ۮ�w
�Q2�ϫ�Y�˷�m$��Fq�Yq�l!��^˴aנ��<���O��pUW���g��
��p���߸�h|���>9Uϸ������cd���,q����zƯ�n��VNE�P�0v���sS�;�i��/����?����A�`+���џRG6���k��a�*�3�:	����@�'_��� ��}J���q#���Q�\���%�h�̯��V��bǀN�!JL@g5�2ہy8�Ƕ�^��&s���T6��	�UH�R������4"��0B�,���A?Tb��~#�7��v�ԉ�z�}�S!X��R���4�6�QO˻�ZW+Ǧ/<[cX�Dm--[>E!��fqK�:w��$��}������e9*�zcgb�13�GgP?^@���' ��+��xP��nc�e��z�װy��鴶F��+�>>O�f�ZaΔ2q�yK��ߗU�)��E�]d���on���0}��W�7 �bXs��~�c}2�k����g�|�*���zp�<6#w�h�o1�>��cP�N�d ��Z�˥��W��`Q�b� 4�J�U�Dћꝏ`�.*���2Bx��}��BG��l�+I(�Rqc��0P�:���3���M,��kL���\l��?��\m�M{���dϨ(P���?UR��Ґ�y�*���T�-���X�E��WhD��PF��Dřݗw6��=�|�*}�hjD�8OE�h{p���_�l�jk�#;	<5 T�_���lE<� -�-����\���$���6��qoݑ+9Z8�(9��K�>ځ���T�f�8�-4�7�\�/�F_C[�81��,8Xg�ޭ���u���:�]����.KȧV�W,)�-ܴEpo�Mc�檑zMK-���m$��9�\z׾W;����`�r�sԇv*±�r<*�9DE��UǬ`}+��di���Y�d/[�̶;Y����:�5G/��҂��t�C���KV������,h�����j���$\h��7Ʊ���T%0�[�D�yƕ�����#��g�&�i��*�]O�q�ڳ�v5����~�^N.�%�n�,>�=əaQ�w�0\�x�?���b\OZ�o�4�)��F��F+�f�s7
�GC&����v氬��l-����j������Y��i��M��8'jN|�F�&9p5e�<��M�ް"��)��=UE�t]��1���O�W�R����i�H~���
��/ݔ�٤-]�7����}Qg��������?�����P2[4m�JZ+/�^��0&��{b��JzZ_�8��'�j��8e���A;�-�H*&�
�*�2�q,B�%x�������	��ƴ<0���ZD��ֵx�H1v]�){"��#�j'�%�5q�T��DO6G�P�
�G�5Z���r�Gmy����s�E�f��i�:����,̆T4M1�Ad���>�%!��1U#C�@o�`W�-�r�K`��U/IQ���IK��y�j�WN��2�/���u�M�ˀ�M~�VT�&���@P��1A�C�h�m�T��pȮ1G�:}J���!uc8ٸ���q��2jy'�,�ט.�=�'��7�3�i�S��94�8������0�npO@�K�?�ȧ��S*i��]7W	�3E�S��0_�f��� �C�^�ޛ�~���6O.E��֥��K	�n��[�l���nˇH3{o��^
�r<��Q9�Q��#�K?IzZ�>�����*<�~�Kpq)@E�.�w#��u-�c�4����,P ��-����I�-�>i����aY�X�J��B@T�~T���������y&>~�B��������VI� ���3���#����h
0VV���M~��m/ˇ$.�V1��Z��	e�Nm��XuK2ZKc��у���/��:b����H�a�#)3�d����y}e+$���	$5@X:�^α3[�s�Q!*�&`����H&DCr�T-;M#�$pa�n�5�`N�����^5�v��!��^�0;k��� R=���k2H�pV7��'���f�Sc'&��(�(�)�@�!�X���͉�q�
M�\(�H�Gz�b}̗����{Q�kˁ<�[�F�b�K^��3F��/�$w!l<HGR���ӏev��ϸ_��������g��'-P@
lw���'�+�A�}�{X`2,T���6��'�y.��?�U7�a������OJ�gn��ʆ��*�"�$�$�G�q�5�l�Ҟ+�2/Pס�J���A�:�8�1�o^�ǳ.?E�R4P�N�@�	 Y��=�F���`����j��p�n��#rzˠ>ˉ_��_�J8�ʔ�#2�����Xy�9�Ռ�6F���bͅ<���n���Z��C�D�k(��&/�v��QmQ�K�S����&�f����0�5�#�͕&�oГό�R0�Ą}#��Cѕ��E�o�{ �W):b����.+XH����lr��_�A�A�6��&4O9�����$v/��:	�ZF��.0�x�������� +��9
>�3���^���N�%l���8p�A��b��MZ���_Z��]8�U�#�V_�e^}",3CT^۵�Lj߃XM��J�� �!��n}�	����Lkc��P������G�셸@Tb�\�M���>���z%lq�:��<Øf�#<M�P�����8p�9��ѹ�+��g���Z�#c�j�=,��m��a<���`������I`�R�4��X=x�R�G�;�4iu��0.
h)��s[�,�_f�,rّ�lOV��YZ�C�}��P\ H���В`��0w��x�c�R^��KuK��,k�~bw�	�)~_�D�����G'�Cn�����q�=�	�4��p�Rj���iH���Ya�G>��xS�TTњ-���yB2�[$�~��@vO㇔��xuֺ�6�s��Q^��Z�˵VЎ%��D֩��(s���&�XXC9�E��W{B�z��-�#�&���� ���Ǭ�.tJwm�q�E�w���U��:Oƺa���D�r��n^gg�̉Ȇ�&X���4����
�-jpۦ���*�@\4��w	�.��p�Ӱ&��0i �tԝ�f��t"�ayz�*�����G UE4�Z��[���"��d�)U-�銱���_G���ug�;��s�YqL���MK�"ɉ�}���C)�%T΄�)=Mq�	4���]�ް�=CL���M�B�&�����nĈ��8�ç>1䀏�v*>h���˱���:3��0��"Hb<�y
_�)H�#��w~�܈uu�/`^��`T'8+���ny�d��G�q�I����������X��N�ZF���a�O�묗J�.�0ؐ��e
M��Jm��p�m�X��l ��I��#���j��]�>��3���{��� �����b�[b94�����`�01C��YK)�V�f�FbA|f8(�ڞ^.�)���D6����Ktm�hx�x{���%�b�`�X>�z����; I��%�{�dPޚ(��R��G)w6�
�#���c&��?HscA�
{E�fج������&�Ų��Xz�����	ԁ�_z�|��z 2z���d2)hd;�b ��ϝ�$8�w./��1�G�w;�P��1�56�e1h'���	c�^N�B%J���kg���?PT�O�d�L�g�
Xwx-T�@W:�m�ѷ�׃���{n�y�!NJy&��g?/2 ^��k]�w{�k�1�su=$�4L@��y'�"���\��}i9qX�K':���J��vi_bg�#$6c���y��rS�n�;���e�%M�������/>�~;2�-ڥiv-v�1'�{�g0g�Df��'�&Ł3�-,�ا ��a�и0{���t��9��������J��I�>\�ρ׼3@��=8�8Ul���}Y�����Bp.�q�mf�I����@���һ�0��RN����@�PL4���]�m�{#�nsg����~!�H+��u��U�,{� �4疋��Ruv	o�&x��
�8��������oIy�0�F-���'�M6@��/��x�m��0L��׮Ǯj7`�ٷ��博+�H�C��9�ϡ��ePǛNxߍ�{'ax �����OޭXBv��7QA���(�3LnR:�<��-�5J!@�*����߬戔U��^}Β��� �
�w>C��0�f�Fpڎ��J��?opSૹ�);ǭ����&@�`K�?K�n*� Z:q9O�n�����H�g	_K�Q$�U���q��6�t�&�k������s�?�iI�	�R�1��2�A4��銟��IOH��G�\�h�k���,	r�nj��Pߞ���ߧ�5C����?���Hɹ��:���B(i3(�,��WV_(᝭����=��^��)��44�� �g��� �9�?҇�#i��9z+m=�u��1+�j�f��kp��K~��9�6�|ƬӞp���;�4[���+��{����[iÎ�Ic��,z��w�^��{����j�-�Z�.�-o$a�aX�)��x,������)�/K��B��F�~_&C�cE�.��^b��Zv�m�[ �U����o��h�+7������p��R)�d���`D$�_q�2�m!���-����.޽��;9�?w��ʋe��J�Y�����<��&x�(d�ˎ��m��Qb�;9P���Wjp����k��$^s3r>x�k��C��zƺ}vZJ�h��O�#q�r_�n�����q�h�������A�l�aQ#To2��HH�-���]s���t��#�p�b��9������|��ɮ>��3�ISP��ӎ)�[\d�A8��[�o��q�C��f��b�����j%�e߽.����ڛ��Kӽ4hz��ݚ����p��,XL��X�C���{nFU�1�������r,Er����~���� *���@ׇQC��[�ј,�[��i�-�Y.v�{�P��c&K�+�SR���q��
=�Kj�.�9�PC�O!�5)��9���a0���&2���#(:苐
8G�D��̩ ��pK4xKg�u�ݞ34U�a�	:���;��'J�9��#"PtN�E��h���8Eu<p��*�FX�˨�)|�ȿh�w[�Ȝp��o�ڋᥬ!)X�}������
��ED[h���O΂|u?ђ$�qNK��J96:�������A����+b7�����ǈ��lO#�BX�n9��9)):�M�9�qf!b5�H�陟�Ҫ'׽�I�ǱE`���t��'���\b�"K�U�V��~Û�œG�B/�<.,���c�Θg�F����I�?ũ�0V��ˤ��ݩiM�Ù�Wҡ�����]e�ϑm�Q]��3�O�:��I�GOBN����]�"a���'��{��\P/�h��.Av��S�V�Oy���ôO0�#r��;:��g��?�`�ҭ���՘1���w�4D[]�D&���=�Yȸ`���PFF��
��q�y�=�	��ɴ:�^W>+!`GBGb�u%�O_��l�ś8���k���of�d�JN����i�a]j�lg4zb+���Q�|�頌�)���� K�y�n��)�O��M�~��!��-rzG�Yk����L>�P�˃��J��n\�%�F�{�2}Mcݺp�D�)�ݕ�:\+�9�+�n�prާ��"�Ŧ���7��`�[�i�F>��~�|�S%��W/�5�v�@ޭ�w='tB�E%8�Wa"����c�ة'N쫣�LtE5��À��@�ڍ�)�<C�{�Jb���ZI�(�@{�J8eu�w�z@����g�6��Hr�H��ݩ@��A��$�,���c��갿q�3p��%��hj�����U��l�F�MMp�xb��^�o�4WJ֫#��Y~����[2�v����f�4#���xM�t�iuH<��{Nb�E�}�#�moҧ��bG���xg���/ڽx���6�PǂW�c:$����p�<��{��W���(E��,YU�lM`��n�l`�gCG�
�g�ǘA�s�]�p���~&�K΂b��#s�]��d��z�������N�xsw�įSˇ���-C���݌�`�I�&Gm����Z[��6ƈ��pK�W��VL�rh/N��$�_JM�i)�k]s���z�SR�"��c���F�t��A]��B��@��^�2({z�Q��t6� �4Ă�(���i�G#�g\�d�S"���x	�.<!���]P�g�gq�k�A�̫Y�����v��yj��Ó~��i0�E2F��G�~��G�t�&Y�jn4�NVbۙ
��L�ܐeJب�����N1/Ѡ7T5d�4t��c��L�Fe2)�w. �p�u.�+�J��)E��^��'Ζ�����j�բ/�Qض9���b*�ք}9!���9��jn`�v�0V���+ �¶��Q�cR�8�<�u� ���n��"'�]g7�E�kbZ�D:�a�xK3�[�pNp�A������rIg�+(C��y�d1���>��%s�P�bړ�5d��Hr�O{g��M39v� �g���Q�/z��Ǿ�v���{i�}�:�����!�9v������S0�EZ/��Z}�����fh���t5x�/pZ���͡���?����+���_�M%����~q)�y�zg$�$�5� M�o�9�� f��(:G�$L�����Bu���պ��Z�S��8�%oFـ[��b��P9  ;1�2�>${�(��.�����h�����3�|Y�6�^�AP�H��9~�@�$��p+�6���tYR�ủ��%io�[J�o	� �f�=��6�5��f������݉rq�ҘY�G��j_{�È��,�o���C��>�sf!{L;��ɦE��)�-�|��-�TJ+�X��z6)�oSXO1���y�D��m!��,P���@��������}:��E]t�m}.b�@�������^d%;��떞���e-�(�����������!�DO�	Xa��I��B���5�.lMC:y2�Te�~�j����Jѽ-�)���D�;�l:�[ lD�p;����?�ӥ3e�*�u��6�P=,�W�����Ε��f��q�?�����$~�h�����D]�$"��/���H�o�ma\�v`����Y�?p�e�Ԓ	C9��R	y�s�;J�D`��, ��4"����ֈ	�� �jGe�?<��O�맴M^�ۺ����p�K���0�3�N��`�Wơ��g@3\-�b���3�o�G�u���7��8!��d��߱vF���nW1���l�3���!
��%�⮷&aa֖��־q<.�kgo�XgH���y;2gz���V�̼K�_ą���b�#!�%�>�(M!ʏ�D��%�A�����i���������U�5"�]�V�����K��;1�|��C�H�������\
� I/~��[�m�8EZ�[\�ז�9��X��*W��!<x�%��k5Ϝ�����b$�H��LNX[Ҷ�,ֱ���kHBǟ���6<ד�x��N �����B��O�	\�X�Qf��F�6Q�j8<ƏG4��7�2,�u#7���$'���E��lZ>q;!�t�f/��z.�*Ԥa�;��Ykh(�Q[�pXw@�s�?����P]�0��/��WS��U�vQ:!�/x6�ǩP����L�:OVݷ4t��ӛ��	
�j��q�����MU2A~�Q�x
5�	넶`�˨�mUxy���(��Ǚ+ށ������`�~'ۚ���o���V(�*��	�D�>���~<i��rpξ8�X_~�8��w�?I؎o���Vܴ�L?���=�C�+�'ML�T\��
R������Ea��}Z�X�I��b�TyV��A��Ȳm(��u����ݯ-��l�K+n�<�ˢ�O$Jy�wH�rC�k.��p�����`���Y:t{s1��%@���m?�ci�Ym3%��Y�U��W�U�7У���Qn�k�� l��X�#���D�ϔ̣�i5��pz6�� �7�C��A�j5*��\+x��dv���O7��'\�P0���]�ֻF�bo�c'��m�y�C�2[{܂
�f�`h[�׍�d+T������o6H��c�>��z�^���N��#?�<�:#���A��� >F�"�����=�@r���M+����QsE78;��G���$�����5Is�[���󈵫�ǖ�7]H��C���Xj �="�X�o���R��>]�����B����A
fP��"~��ҞØ���,g��7aJ��}1�g��I�f����v��I3����d�5��@�#�!��-��(�2XCN�&F�0�	ӏU.��?��C3lg7>���me˻}�b�����%C���=�Q[!�u��2]|e�,ڼ�/�R��bl���J���9."g�˹�1�X�M2�R8~�c}~ǂ ��wς~]Ot��RTu6|�Ĕ:ϝ�g��y�g���� k��0�+f���Pnm����o����ɺ��eW$���A�#1}��.��c8��@�>�^�\���B�9i����R�V�<�N����CM:�~�@�t��,��EczJ�����6�����3� t�C^��e�8̈����%v&ma�,�,��P�"O��Mx�>��Jd�$�  �=p��4�����s�҉��W��i�~� Qj��q>+�n�&���c�
]Z�\���_�?�;�?NU��hJ���WM:o�Ki�Q99�^T�O6��+Q�j�ᗔ�4��wxd�;�������ӛA�m��isk*�]��s%�Y\X�q5)�?�͋VÎ�o@a��X���x#[�5i�1xs��� �!�J=}�hdO�����1��}���=HH��<�Mv3�#)>�P��V��@fKȺs�j���r����#��?�_�`��'VR�u�E�8�Oo�q���ffV<�Ґ���Z�)����q̀�[�S~1�q2�!b���9ҁ~L�W)����[d��`�v
�L�dd�n��zY�b�U��h��h�I���,�9c3��x@�>V6�L��p�׹g�)�_$^MY�x��鬆����a܎  ��^���4.��%����q?�x��8��{�F���k�l�8
+����!A�%�R��X61�J/!EF�-l���UK7��#��A�d+��p�~�BT\��t�H]\�7�;����n���xk!.k�"<�z$#�����s�����U���}��F X���Q����t�e黍`��N���1/޲�l@����G�.�l�bM��h��"���pՙ�H�'5�A�V����r4��_}�"}ж��?k���#�A^��TM�Wsw��o�q��+�>�^�u�1��W���I%.��0��B��͂��&���jW2a��ƟG��Wn�C��ҁk�;���������d��\5M�<����y��� s�X����o[O���
��^���	�`>��+��22�F#�t�Y=�S0VK�=-����f0����ΈQ���YT�oZ�2wS0�=��B
�̯���2Q,��9/RfU�a�h��0@ 0�M�� ("��֊>!���Gj�O��qB�I:���d&Xa;S��+�������s	tN�]ME�G���[���6D%��O�6?&�5���ӫ��d��Tޟ����[��a�� ��4��;��zӫ��yTQe���J��*C�G� =�Dۢ�Wz�|�@�2�Б�`�q�e�� ��?�Xbן��2e���^�]�`vk`�C��*{��r(@��}	m��w��/ 	���#�����ΤQ��+���\� ��*XAg��y���������L��B�.+�CR�w�;�	S�Z��6��D��*��L�qﳳ����c�\VS��F�q_�~ڐ�D޽A�-�����HN�����v����|M�k0����XL�ѭ�b\�w���3 ��')�~�M0w���|3����U�U�9m�D�����S<�B�6C ;�u�=��bc�u���)�B������u�<�D�gw*ҋ
4�d�A��{TՊr�L��{X˔���16��/^����3��O�� $�2U���\�@�?(;���G+�euM��* ����Z���g�����y��6�0�֎Lj�gX ��;����ә-|�N�u�^+l��E9R'��4J̑L��j�Ǖ����W��S�}�[��M���"_�Ot��]�I��➻i/���dWȶ$�`
��>.�B)����-��>ӓ[���ڐ����r�qNcY�ϣ���F�a�}I���y�4-ތ?�f=aY/�xM;�8��݁	nu�J���{;�1�;�T���I^�o�N����?)>fG~�#&ɜ���ޖ3�^j��>?!"�!lΌU��(�<�m�^�ǒ��c� ��>敂P�Z��Ժeˢa��y���2)7�� ���Y݇�C2�K��k��a�W���	b�w��cr��i�˥��Cy.�qh�sl*��ε�+>�T
]-���Z{����Ϸ�!ʵ���X�I-0� �b�Y��1ِ�MV>Fa��2z�s��5,w&fdNk[�u3�Z���^}�/��K�&������n#4���HI�5(��4|Le둫$�v�Zx�}=޻04��}���ٱT��ܶ0�I!`6u$�CcJ���r@v"a�f��v�cI�4J�	3���#���z��3����ā�H5�	���B��_]�����Q�9tL��ᥩ-y�INo�I���X����1�ѡ<���7κc��g�_ҵXN�)���(�tLGoI���޹�Uو)xO��V���ƃ@t~ЇR��7����Nk����a�D�L5k ��m�������Qn�����ߔςc����q|����,3Y�!� �5т�|d���֛�D�}�Х�����X\�(=�������U��YgoRG�-��'F��L�����=�fp��_c�l\Һ��ϕ�k��h�hv�o�	_[������à)L��\���v�r,��/�!�k0Co{�E@��ϖ��(�p8�� |��z�.�����ˊ��� ��iK��/��zL��0�.���_�[そ�3���W2��)f�~:�E����x4.'@��i�A!��0�~ +W�L	�nT}�'��������wsB}=����]�Lm����o7d�5�2>���?�(� /�zr�{}p��4���|m��ײDg�bV�`k ������	�c���&6`�}n��b WN� h%C��}�k8:p<�>{���8�H��J��sr�