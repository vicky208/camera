��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:���[�S�Z�7����*�a?��%8��Y�a�z ���P,�lN�/�/�߀ړi{�,ب�ɬ$]��Y�#��J'Q�D���^�ǆK��_,�k���Bԃ��P����P��������8�0�@_\\`L�2�V~,��h#����[��/\R)�8e���VJ��ҋ��eSǑ
���&�K
����' ����tg�%0@���'��n$p]�b]s�3vM���_�~_����<����}Sk�[���g��B r� O�\�^�p��4Љ�����Sl�m>��K3x�X�!�fc`bKA�j	��8	��Kh_�ݲj���/!�D1�����ӱ0���〬�[!��)COr�~ōg]+(�/dR�0S���2T�1ĩ��y?�cPF�Z�9z#��X��CZ3�ae
A�l3a.�H����H1��r}+�C�S<C�,p_��\���&��dH:{3-�
ػ, ̭?��?7��+�1y&m�S;2�fl�4KcKآ��\�2�+e��y+U���<�|�pn�Oˊ���y��+Xe����`�}��]�1P��奭Ճ��(ƍ�@�Z�v�>�>lp?���Q�_�mi���Jz_��9+p��o���0��r.Po#96fF(L�,X�"�AA�l3c�w�4t���@�j���q��XS[������G��@���9�	R��,�*?/�n�s���e�����)}C�JF�
��N�R�I�ԏ*�õ�~��
���1�`�@��&U�[���M��	�(�k�>��b��3?��gV�6���<7�t-{>)��?�n ������}|9h�q�1>/*�-񤛤����tƭ��JхY.�{���fhރ��v���_�M�"��S��xGT_���u��Rr��O���X1!Q"׫�]�O^�LW�}a�l�T����ev��/�2���w#j^����D�2�7~Àn�VuBq�㷨{Gѝֹ3R�F���9N��n]��������'$��gY3��4k��dD(E
9�zcx�WU����}��&BG��U`%C�Ԛ�iv25*��F ���? �����۬4�Ń��X�W�當���C��pl2�_	��*�x�<�6�f;+�j'%�-49к|�ѷ�=�f�V��	�،�[���&i<Wf�t5�p�����ʄ����HY�=:�&o�7��S��Y��9��j^�����Ju~���@YCT�n�ţ��H�U;��~�!�j0�ʎ��ݺ!�8�sVU�4xU=�m>�V�9�E��D�t��3��v��z�f���;�/�M{�ݟ�<�Ye�էT��Y������cJU�;l�cP׳l�W�e��^��r�뒃�k7O|G��2x�9��H:��?���W���w��#n�E���>���_�u;��ӿ�471L��E��������;Ağ&/a��E�Vv�,�ۮ�q��n�p*���?{Z���Sr,ॣ�#����bеTYo�M/�M�;.7��P٩�oR(���I���L9:�No�����=lca;��RS6��-Őe�!��	D}���[���
t;����g�4Y�jDVm�n	�`��Z1W��yZO�xPhK.:pPb�O;G[?�6_�c��H��?�ƀ�Q�W��N�ڤ���a��F{�c?�3�[ou�,"{���w	 s'QV�;roeB�+(��z���Mˤ���x5Ox�Xr"e�����/�H�0�EM�V�'n�@渏͹�qq?:�(�����p����s��S��^\�"�c�E�A��vw�[[K�
�z�z�d
`v6��@�]둼d:y��ҵ)|,�Fh��h���Dr����"�N��c�YxW�ˍV��O&%k����O��8Ykh*YH�(5Lߵ8�^�]�����7�xɖL�z�U,
!�U��ai�1	��=��� �c5�g����B3� �.&~Z�Ú<��8�z�!X�/B�a=^!��?2XX��+���)�T5[���M�;3n�@�Ϡ�m�R-�����_�����9�����
 5}w} ��"�B�禮�U��~��֩LcZ.�Z�����A�4����E.7�O'w���,�J?��h5��}�"���D���j"��Ta�rZ_�7+A$�Z���ȻF�J	�-����i3��%H9m���;�4xN$l�Lu]}T�i7�p��𪣾ɱ��J�)��ᨆ�̋���`ů�Xh'��\5FE���!�[�ǘB�9�¦�����cN���γ!�&_�^��8���7�#�-�}��.��t�՟'�R����U|��þ�^5��<�{��:�g� 9��!^�3��&��zJʀ����o&}��t�٥I�n�9z�Ғ��%�p��{�&�X1s<�n���#�E󂬯��aߛA���M��hHo�=��lu�ZR�����I'�4oJ9�a�м����>x4z�Rf���ט9+�|� Z��� ����sb��Q6�� x�S5���y �l$�+j{/iK58�L�Ԯ�>e(�w�
@��
/��:"���c�en�i��+�RG=�F�6{���Q��2�*M\��OH���H��Cr�/γ�.Q�T+���3�7bx:����q�! ��\��ǰ*�����%Z�P��5I�HJ.l�˜�}�(����������p��EF�6�b�]~g�S����c��^熛l�2�� I����{�A9k\W�g��;ƴL2����>{���-V���%gg;l:�+��P]��`��N#n��(=�O�U~9_JS�}㷨/jL�f�R�|����x�0�q�}�qzo �gc��oc�%�����os���1pc-e��?����K����~\�T��!��8�bA<g���ߋp��\���p�8W+[��gu�N۰��� U/7Z���W`ڑXݣ[�����upͬsgFA��a9���L��g�|��.\u",���'�u��sõ. �.(�$[@D�7��VY=���[b�����u��(��>I����}�@ �SaQRw�R/,�.i��)X�/n���'^c�b� ���^�+��)Զ�q����Dgs���=��j_w����kt��9�%����������/�'�RCF�����"�VC�%��><�{Y��@���� �*t�q�u<[��RCz:a)�_[ѵpx�)%�|�f�Q�q�H.�H��oqЊ�K��s�����@��a�b�l��#���p.�w
�/�t�zd����ҷ��J��}��~����VW�}�O�܌�:�v>W�z����'�z���q �k)gV�0q��[�ԨTug��S��q*1+�,�{���#�:�Cb�mեos����
=��	6��^I��h��HKgl�G�;��f>L�:o���p��x&��b�$��
��}�8~�t�D�`G��������G-c�� h��cC�,W+%Y<>��t��e^�}��&xÿw�eb3�ӧ����]+h�X���?|�6?�v�t��DF�F���S++o�aUE=���*��F��
���dIPBZ������{Li���%��c�/��ȫ��n��gKu�N��ו��.�B4ų��#h�B�t���($M^�KIl�O/OG������r�X�}�||��Tw�L�+�QO3�K�qN������)~�=�S��S�dvJ� ��|D�:�-ڼ��wJ+�E��5T�-a�|>�JNn����i�_ N��!n�����q��=���	䚧��W9O�w��,�Gc�u�e
����S58����&OU��k[��(�u鲇#�ALm��`.� A��I+A�7˾th�j���{X
�n��������T��iLs�~��W�/�Z�55���,��FپVbFr��]�]?�?P�|�&f�Yqo�F����=��-�c��i�6���W\9#9��SZH#���!��Q�.s�?�E����3y���`{�h�Ŗ<F�\g�G��9�o���%c���������\�5h���l��T{m+�.6���6'l��W������Y���e���2v�цr�8'����ʨ�|�O&�險���e�r��pn������Ղ��=l��+*�ˌ�\2�s_�sj�o ť�����<Q��塼���4{0�zc�)Ԙe���Rc��-C���L�"���-ՌW_؀(�3�W���w2OpKc\(~�ʠ=���f�	�t��!xM)X)�%�2�t؃"RV�à��X��%Nl��!�EKZd�c�P���~���y�~Ɨ0���XHA��ǻ�z!��{�b�C�A;� w��cs�a�	���>�����"�vG &P���Z��*����3����y>a�U\O4{�0��PO<$A�!���Ɠ0h�wZ��BG^�'d���hؙ��<H�)�P|J�w'�ua�v��P\�T��.�Dn�<{|'0��+I�j#-6�W+�b~I%#](p5�5/�_�F��VN�]�����&��	�Mg Z��PT�_�+-CJu�%��b���G��lY�Y霺�?���2E���������#v�C�O�@+���p��]�RUQ���"֜�<ac���_c��قS�O'JǨ6���ͥ]��6�,�nrI�_���ٚ#n>ӟB��<�΁l�Xk6��fȼ�SN"��:���Z-*��qp�V�5����FGs�[��!n[Պ�P��:�l*�l�~-\�����*�����6}�kG-A����r�+������"�o�d&�礶�U����*:{c���`f|Yb�Kr�,|'Ŏc�9(M���(���!���c����Qe2.��mr�11'�CՀ��0�&�t���g$��|�Y�V"��Ӭ��A_�w���衸��y[�nI���{��0��M��R<�Xω2!���8�= ��?��a���=�L�'ݎ躷�@[�#	#MKx��w;Q��:���<v���~����I	����#w�U��M�U��C�E��-�Ӵ�9��R'
�%K��r*���$Y�OIF�\�=�R��q.�[Mco�vHH��$r0�%�i�TJy+�M�Xz�&�¾'}�K���eGȅv�Ԕ��E��ڵ`;�Y��l,B,y7o��Gv��c� �`�]��t^ ��j	x�$"O�~�Z9�:|�����R���m�:v�y�g�/�ea�ܚ�$+h�����7%v�2BȰz��Jr��" n��ϑET��/?�����~˕�a���\�|f`.�絾���j3 �� ���c]���.���u��5Z�y-!cK�\�p�B<%���dH� d?�Qk"r��p�t�G	�?�T5ǎu	���[���1+�tY����9�b�kR�t7��_�IC@�����:�8�
(�Q{FD�����F���#�G�H�h	��|(�o����g)����K�8�C��w�3ēLà��#��h�0l�� k� �
��2kQ��>%��{i�^�kLT֘���We�)����P����=�a�^J�I/���XZ�������Q�{kCb�1�+#*h��ؒ��@�q?|������RY2�x=:���U�@����������\�oa�*���.�rzON�^BC#���>���r�W�U|9�Us�]1P߾�P47�)��p�ѦՈ���4�/�rǣ8Lc��JhL# ,Җ?������.�V��f\�Z,��g�+�d���P�+�!�=�<Zsk�w^�+�{����j;�H����jN��r0
���� ������oR��^��d�$��;�dI�'̬�TGX�&��J�Ye@$s�Х�����qn�����tQz��:���&Z�z�K�	�M�r�:��M�c��=/5fU���c��#yf��*�Ǧ�� ��cᑖn��%�� ���1Z8��h���v}�z��7LCF��H��eP6�ߥ��OUjT��p&�(n~Zu��|T�� �L�1 ��M���|h��9�Ca:�����p�ۤ��I�l��(�ҩ����qhA���E��j�&�?���l�n��M�l��>�R��聚y�Kn��c�P_�R��tWÒtLtk8�1���-ç~{O�d �ѧ�6�5�P۳�VJ�싿���^�a��5l�he!�"a���T��,qև�d�����bD|�<�, �eJ\�2�,v�H��s��=���(�:�^m�c�( o��z�D$r�}�t�;Q�d��k� l��D�����UƪA���AN0����ltDxwF��5�4�+����T�~{���h齳��|98���PQ#����xrt�O��d��]f���*> ���l{u���?m<���M�RzYބ����5�o��ӹQ_>��磏����ѕ�<C�>�楼�i1��_��-''r9�pL4�K�\<|�W�&�v{��\6��.�2F�'Gh�	�d.��v���E��؝�i�h�J�$��OIIx��~F�?��Xm�g?P��U��4��v�r-�H���G��t|- �zv�f����X��
&�Ѓ�rR��Gd�Ba���$�ƈ���gUP������-B���7(C5M��S���@�^��Yf	��w��<oΰ*_�y��=��E}3�V g��pq;1��y�~�Y�Z����s��E4z��q)�@�&}��B�%9��R0M��\�+c�xKi�f҇��2e���H�|��\k�5U�/~H>������Lr��b��bX�a��ӂ�$�&�_�Z�%~N�DJ�lͻ)~�����r�&,{W��5�g2��q.��K��_��}Mqy��.�ܧ�6E}-�ѐ�E�9v{���+.�uF� ��L�Ny \�_=)aI�\��,�-ڹ����2hvVe�|m:� �s�m��DF�>h�G�(N�q�AE�>����R��,��xb�asJ�,�%���¡<�EԖ�x�������ЩG o(Β�3�C��K@K��fQ�x
	��t#}2��	����Y��oJS��b
=<ɔ��^�.uL}�p�г�Bt���ԏ��f�3� ����-kF�)z����1{�*s��0�e����Ґ�we��笆d�����HD�j��?��&�;D��u�Y��� <�+�W~B��/М2��(��� v��n���K�{Q!�#m{�E�����7��������U����ueDXR*��H�R�bl+R,*�Q�\Y�&M�+{N$]�*�:r�ۉҠ���JjVʾ�[��KJ��g��L5IKv�::b�`6��bV�T���^�;Zn���B�2�)�B/$��w����@t�3��p3��]��@Ph����R.
�ƙH�({G��鍧��8�J�|dF]�x���r��So��q8�����;]�f�e�i��i��v��8�h�S-n:->��#�U�c�r���c��e�a��v��&�,��g^�L��Q�͗S�^R�����$�a��Wl�qʆ���
k1�tBt�1x�h}ҩ�*�+�U���&�Jx�6r�e$��8�k�N1�{L��.�嘼���@��u�@*7�������Z(E���i�ʂե��6���Bq(�d�EM���(�Tn� ��H}u�|��.?fu7I�����h�n{]3�/�8�`�> �m�0��,�Mˮ1��ܷp2J�V��Nm�ivi�ش���Y��$J���ާ��SK�B���-�����HM�'��Ty.��/��L��ޫW�f��rXV `6�.=��I�+Nɟ|�`B,Ft�"��bHaG�"bO�Ќ�d��E;�E�ք�������kA#�{m��Q
E� �x(J���+��� �[t����������w��[H��F������1��UˊDz��7�5�������T���&����'��Ӂ��M �/�߆O��s^F�YJf�&��}�Ղ��CE�g�g.�'׉�G͡�WdU>���R��Q} &T��ҷ5l����$L�7�g�Y�5)��r
9ʀe�����9�!>Q���C\'*:��A_>]1�R�׍`�'\Μ�3㋣̠�h��д�?K8K�
�Oy!�[V(�{���t�� ��`�"#��{���|�X;Fb^�m��Y���l�U�c�x�OV����?G�}ai+��������h���N`�*W+Y/��ӂF0%w�8�QO�U�?\��Y�]AZ�.	�K�:�;!����l�������^�WE����_��`HR�����o�ꅾ<*"T0�T����[����`���t����d���^�i+�؏�g3�L����p����\��L3f�q�8��a��Bd"���.�b�-�-q���y\f]0��I�-K�k��6+Su�g�=���6r����=�M�?+H��R�9P$�]�% ��`^�ca"��X�ko�
�{a����	�|d/F��5���[.�Cy޺;�Y��2��`ZY	wF��.��p�܌���P�W͉1��X�0����P��&g0�BV�����^b��ot���|���z <y:�i�W8��v�۳�!�"#�B��n��!p�g���1�e\�_2c���c�ƋL���Q�p+0�Oqo����w���8g��i��)\��K�j�Ꮼ�W	��0�� E��p�Y�F��qu�$	��JN��Peۂ)x���KL��(f-8�/C\��r�'�	8�K'E�.y�|N��ش�t�>|�q�=����_�����6�܉�&��d�޸�T���Q���+H��]�;P0L�	X�X��,�`���:��T���{�A[��M�2��P.��q�q��F|^��N��*��F�<�,�˷�����8F����\JL������&��z�+[W�,a�9T�}s���C���|}���r�\ͪ���̂���.QM,�Mik���ǰ(��܄X0��ƴ<}�M8�_LYe��)�K�V��B�ҳL`�z��a�IQ%�8�i^f�U`�,����M���*��Go�O>ﻇ?�TQ>�C*S��[�3/�
���|����l�_���jOOYi�[3�O��A�Ǳ\V^{���~������,�6z9�c��uI�h��?��`:������w�s��-�-���H��9���f�?�F��g�?q"��=q-L��{Z�Jj_ L�"��π<&kO�"bXH}��>ur��{~Ӎ3�Y3b�m�M�Q�ˆ"�`�q�=𶸀r�V�{C�P����4� v��2M
���X�C%�C5w�	d۟���1z��Ml)��i�&�GF���C�Գ�!�۱/�
��,��9Nh�t�ڄ�e���}R��'4/��RÛ���~�+le�U�.�h?������mt�O�[�l�:�`��8r�ڣ�����s�Xf�Qo��2S&�{$fƆ��Ԑ��x8�*'y@�x������GF��1G���+ ��}��Y���-�mJ�k�.��mo��*���V�+�"r�3$#Sm��a3���oA��n��8i��F�,��*��)�9,~�LJt��բU�$T?D�1�Y��[��B�r]wJ��o������k��H�L��"��X��4�T��݊��F�ʶ�{�5��J,�ޞ�?�t�)�/�9*K6H�^�	cC��Qe�e�����`"���i�¹�[~Cf9U�dD�U��V%%�ƣ�P�B5�bWRG�u"'����d�ᩱƤ����W9������%EE��{���U��D7?ӹ���#���{ [ ��d$��/�l�6X%�N�Y��b]�ǖd� �\㩬y{��Km�}�5	Z��ȏ���fZ�T��놅� ת�����^b�F�4�{� ��x����y�aH��AI-�r�L�\�1����R�:�Y��N��DC�,�a4��G8�ѱ��Wh��[�|��A5����o9����O���)���{_;pQa�>c��ij�OZ,V<������a�)���yF�ի:]�w��<:�Oh�F�R�7�Z�Bf��0���V��Ư�����rj�"k�J푎���=kM��4�d� ~zt"+�~HS;�L�qo�@���L���3���c�rM�!fл�E���Ym�����%L�����Խ:�'��@��H�:�;2~y���/��V1i�L���3�p��uޚ������>��GF_�W���ùAj�����	4�mN�諳sg�`7,� �!��G�و��Ж��$�â���&eHt�NXcN��C��*�E��k�j��G��,ZZ'K=,z����a9�):y?|h�]d0��ţ	"V��i*N��/^��l=.PaI�r�����PV�mz���{Z�`�/��>r�<����
�b��<��Xq8�z	�o�Œ_�W;����]��|=�u���|Dw�O`�,�����iߡ��X��r�&?�A��6����&���)��̌����(��t�Ǆ��,���b��Ì����Mp�����Jo���,�ĥ&�܂Lc�؍��:�	���"P^W�e.�MX�7��"~��M�[���<�m����S]6,$���q�_��~%�>���NXs1't|�a6"ѣ��;"�$"�!��0��<Ӵ�ߨ�>]^dR ��d�(�&�͖}�;G������F3I���z�k��o�#+���e���Isi~����+��+f~�m���8��F�K��n+<�L�iR�ѩD8`YA����C��W�$�2��)��)�q��3���k�Z��V��Tޘg6��F�?���E��2Y�����a��;��'�_v"1g;�+V����_(�&eB�AE�8/rkS�9=Ɉ�uN�����5�r�jlA���8-����+��o!�C����P/�H��l&I�칷�F��:��J�x�q��Z�j��R�P�(h����0�~U9�	�4 �O�~h�o{ս�F��li[~z�'S�vʓ(I.��������^�0]A}� �!i�XJ��}�|�	^
ƭ�O��Ǩ���5�ROv���v8���U�(L���P�����	x��Eġ'��GU��+����Π~�=�B��Ѡ��q*uy�¹,Z�2�$�I�N=)��#a/U�.HKQ?r�4���Z�	x�t>�M�%��N���FbtE���o7��u�p�q�.%����EH�*�.�j� �E����P	���ͩ���D�4QH%�;��O�0�%L�G3��cs����<q�����w'�2����/vS&�T������P@ <Ոx!�2�~��E����T���1ُ}��e_}ՊE���@hC�67E&��'w���u��\f��O�cP�8ߪJ�ɬ�;</=��b��Q6Eә[W b�tu*�� ����r���A����;@(H�s���g���Yn|�x�Gt2ӌ�7�j�JI8���B��b�xt^;f�7~9�{�F绮�+������V�`c����=cdG 5��˫lBI�?�TC_����!n�ouR�@���Z<G���ᤗ%����Z�Z�+������z���E���)��%H�/�����	J�4����P�Iy`i��q�Ö�+�j�;c/��	�bv�9-WU�?��-G���/�O�C�*���V~�˹4����n<n�)�瞙��1p
)'�hqUA/P��J����Ri��Y��5@�0v���5�
��Ǉk���y��P�?H�e�p�Q��m	��x۶`|�`���t���s���`ɩճ(�S[�/s`��Dtk��	�U���8�8�w��Z�&�ހ�5m-	���xi99|fM2j��D��R�-��f	�C#�Nl�5��j��f�fwaz��$���၅:릶A�#��9�����A�|���w�Z:Q ��2� M�,c�4܎˭�MLj��a3�ܼҸ�VR�qSi�E�����`d����c���,�R�{��X��o�?���iPz;�l6�M�Z�z^_\brm����b�?8��icj:��Ǐg������Q�eV�>̺����G��&�>v�K�c�I�!_��їܮ9T�+� ��ņSH����d[*�|�c0k�`X&xI��P�� [���q��gw曣Kx���˙��Y힠��H��&2w���z�i��HB�)��s������L�t�{�S���}��BcQ3�s�m̭D���DnSY����q:��
��5���9{�&ʋ�3X�m��׶C������<i6i*3k/�0dV#��>��U3�[�Cª���҅2�p?��Bqf4ʘ�ET�$��q� CO1��v�!�j��IP�0Q����o�;QԀ�|�<#'f��v�1��}�c(�N�}���~:ɤ�o�F���q�AW���1~�Ygj]H���u���{!�ڼ�1�v�A!��0r�ݕ4_<ݽ�ޔ���9�+WX��x�7���_�Q��Lt|����:���68���v���>��!��T+��Ɖ�����P�t�=�F��6	��&M)g�5��g��y�+�B ;��/�1�xQ]wg2I���x�zb{�ۆ�.M���̶<���T+f��׺�W�i��k�F09�=[2�{N
k8	%��X���g�r�6ҵ��s��3��O�>�C��I
@%}7��
��f�hע�k0�L;tC o49����cQ��~�����]��kYzPw��q��u�IҎ�;&G����������N�q:⌻�߇↮�T5K\'쨳Z�2�����Y��P��׾�T |���=���&�P��#��w�Q"�G���w'�^�46d�Կ6FO�4��r6Տ+��AUNҹ�ڠf��+[�WOi��E��e�⟕�<� c���I��2��W�o<�x����w�j�n����b�3�
1��:u��@��Xr�$�!Һm刏b�]阁�?Ϧ�m��-��a���9����R�)������[�y�8������}{m#$8��G@�c��!�k�H�R�
e<ȳaު�P�.r)�O|��گ������x��o�)d@������U�x��C�D����U؁���0rn~Q|�m�~������s�m8P�T�.1�`��8�����g��n�<��3��\|��BM�� v��Z�⌳�Ic /I�?��U#$g�\�]�����
�!�T��Z����~�WX�� "5����K��mD���\��D�a'{��L˥�2�Dv��r���+�%� ��Y��{iܫN�P^*}t0a[����:��w�#1�Q������dm8{v��v�4dȳ�~�q'���<�v��B =�B>9Vè0�D��ɚѭX�d�ME��iA�D�X@W�I��|�t�|ߕ�GK��)ĕ�;ٸ���vV�y �Im�l�����u`göjZ=&��QN��V��a�����.��C������|?7׈c-��F���k��*�iL�@� ��M�{���A��,�S���]�)��K�;�ۈc}I�9^S^��ypq���X1���xt���X�dT������k"۶��S���'��t�?�,f��i-��g�{;�Ϋ�t����d��Z����IЇjW栬�hq�e��=mӺ7�*�/̺�~�`��s�qW����Ҵ���׆��i��)&�& �Ь�V��7���H �6V�?�V2�Vwn�,v��wpf�]�!/PD�=�_4����g8ӛb�p.����p!t��V���E��=)���[�)x���$
�7rW��;c�����n���Xڙ�;QD���9��@iM�m+*r�Bg�DO��b{�'���}�wy��dlp�J'a�����G��2(�3����\N�k�{�L�\њ�A4Z:��gX�	�3�������ϔ�Yn/��.�!ȥ_��F���-�p�ȅ����S7cs·iFM8�|iaF�{�`���.�μ�l�PN���#��s<~�c�`:���-:�����';���.�/���"V�)��IHu?����m;�ഊ=͡\3��[���"@��/�1�A&C������/f���ru��ʡ������9��Բ��: �����e�n�=��	s,5�Х|�`��I��u�uo+^bL�\��T���x���|3���}x<sܓ���PK�ۄ&
�jbf5@�Ł��Ōf����eΙ�g�{4�r^<�����٥>. �[�i��F�"���h�k'3W�,f]R��X+)0Ç7X9�
N6�������CEpqc7��;"
�q�)���.T��7��_B ]8L��"�K������}Yӏ���8�b�w1j�ki&���m�m��S�Y���LS�j+
b?
�,
�k�Ц�Q�b�-|A��D���c����Z^4���uԿ?PC:`�j�Wg���ַ�	ꊔ*��G�MS
0�CQ:FHJ(	���G���m���-�+�E{o^-�V$�s�S�U��:��+�E/%�>R����\�;x�b��6�	���AND�m��H�3�v�t=��&\��\�@$�'��#��5�a=c��2�� �Y�2��K�z*�<	 ��(����ʎp}
xS����F2��D��d6f�Ҫ�Qs�J]k�z�۵M9!,���H������1�-!��g�JM��`5�J@�j�6���U�fc�t�T1`f��v7~~��2��-�tv�����R #�o��7�P�$/;�|�unTm��)B-�V��>��Vq�rf�)cM �	v�Jc����Rq��>��!�q"���H��*A���rS�7��9��	]X���[��:����VZF���w|��6叭^q3�ǋ��/Dl �k�d=����j������&��{O\���b���(i��I�~�!B"lBq�#��>4<N�u���U�O����oZ=���;ա5Q��&������zf�k��%��zҠ�|}��qH�}�.�{�
7�F�.�i��7���o�����G���^�~���@dÇk9�����[7��|�8�C��_.]�4�e�]G!�ό(2! ц��:W�����?���b_#�"(�]����P�W�?���>�j�P���׵�J�}�)Ö���
gR;���'<�H}�<���õ�A���G���Q!��H�]eï�0%�����yv;�a���l��M��t��md��s�����&̜��¹.��S�!%=��u�3r�A7_��/ٖe�JuO��ȯ;�J:Β�i���F(?�����</OEQ�Y+悬��k�@`8���d��cI��EVy}��ϊ0�S%7�1=1�G�޳� ��Gu��p��""|�(�C*�����D[��ZB���҉��-�U�!`�yp�둊��JV���m��+�㳚��u����᳧!�u7��Ԩ;hI9��}�s읗��r_Y��G2����B��I��;b:��9��HS�@���^ByY�}"i��X���"���X3iH��CL/�
E���)�14�t>�e
������*�C����Tߊ�;�H���9���K��yy���^ylբ���4/�BG����A7?M���V�{.=p�����[�����~Q��5�Y/�`W�ud��y���#�Z_��Ţ�&���A'A5�	ؾ� 7P^�7�w[�k]V�����#o�
)k���`Kd��e(����rT��t�AC����-u��>~�"�j}´m	���=�:�l�+yO-�)}�`��!���բ�� L5�k9�q�R�"��l�"o�$+p��?k��iU�m�=���Ip�BW��@�ctb�kZ���.'�}4&w/�M�{�qg�m��ثؚW��J_�Ƒ%���h�Q���'x�N�
��0�t(
�z�(�םܮ-?A��$�ƕw�S(s�1�<I/E����d��I���U�FQŀ����)�8'6�f� �<��!8m ��V�χ?){��L��� �&1c�6��R����j��-�ҋ�f/�SS/^�D��-��[��S!lo�ƫK�-������/��Do��Ǝ*�ǆ��`jS	͉^D٢8J"����~*d=P�I&Ĥo�@	�?��=��������G�Ҩds���yF� �Ϻ������#1X��ə<���,kݭ{tNq�����(�#~-�=�L�(����p�۰͋��-+��g����^�dF]� &S�(��B |CA8���!��������;��Y�[�.:�dɣn�_�#,�Pu��݀6/�5�8cp����\>Wh^RM蕵����w{�<�zN��]f� �9WF�P㳙J뿍V���R(O�q�^��j19J�֢����Of���2�e:����M7��y�O�q���IXY�I���v~�X�Aj�L��Q��b1��zP#���F�%0�2'���$9հwo�}OPw�"����{�'e�3��RŰ:5g�W��͊fN�K�F����_Ap�!h��-��%��|5�l��[��m �{Q�3	���<)<fi��Y���K\\�C��2�HgS�kB�dL��3��,UqK�.+�ڃd��\b�����??F��6�z�@�EnKɚL��0̀܉��h�}���ɘ�ί�9qZ�.�DJ(��-�xו ($�ĳ��=l�ʹ
��&rhf�5�Ku��K;��+�Aۑ�X�l��>�^ ������^�fX�B(a3 ��g�-���o��F�=�)^ha�iT)�c��9���F��0�q�S��|)�c�.yK��t��/A,0�]@Z8=��!H�ǎ.<w���Eֹ�w����pױ�($�Q��ՄP�ݢ��Y��;)�*�r�AI�)���H����V��w�us�W�#�����Ɣ�9��c�� |�����2T|�0�������\�n{L�����;��� I6�̎����}�K/b0u`�jm~�W���鮾��4S��	ҜY�ស K���$�dZ~�O�ťuk(��X;���/�3��㉫��m'Ȋ�;��8�G���y��W�6�a{i�� ��!V��K�/��Z!vQ�.r�H�Q�G��cv��}��wʳ#B]Be�U�k�mu�����[3���k�;�8�Ƶ�V���̚��`o����R�k�����(d@D��L*�Ԁ�+��t�����S�Z�/�y�1S�O�q��Տt��K�
�Dy�8����&C�䵘���������@=��s?g�N���7ƿV��YWq��xXi^�o3eG��4���뾡�� ��jW?�!��[ձ��Y�z���6�L�ĹGO>t&����	s�p&@�����đW�:^��8 +�$R�_F+5z�Fp��vdw�s$�	<��B�m��~h0�������q��*�=L	z�p�����t��y����0�3w0���5�!���w�q�5������ft�gQu$
x���t����8Nw�
��:��S�Ww�p�pkg��̒K�9c+��s�O�Gy���S�a��t�&+���<6�Ú�Ξ�|�M���;����8�X"����Ao����s��L=s��,�?�[h�=Ҭ9�G���mƕψ���eS�A���E@�̵M��po:�>"E���r-+����H���k9�c0Ę?X��=ل����f��tZ�H�Y�i���+5��O�S����5�м.�g�yq'��@!"<�h&��{��τ�Mu{���W[�îFhܙ<�Q��|��>ݠ!�xpy��������O/���q���t@��)��f�1t��5d51������a�#T���PW_|�{Z,Bz����
H�ur�����9 �Q��K|fJ�{�@u��|�������4���}[tq��59�|
����4F�F�J��h�jG���U��PP����_�����.eH�c�(O�"S�YOlQ��b�v{̛p���1��yY���\�$z�n磑/W��6U�P6�*$w�q�/Pמ���u6���VO�ك|�K�g�z;���Nr6�������e\A���鹭q�2�}��ф�vL��A�%��1Ք	Mܯ��`�I>��
����9񝻃�U���[�F����n� OE
���V�����cM�`|k� F���I3(�,b�������.���Q�7U���P-����Q5�wKV�Q*y����sV�u���݈<3�6����҇�J�:Y/,���G���8-;}�:�Px�iӖ$�3��
%1��-�,v�l�=�pC���;��\��1JjOX�3��}�y?�LF�"����	u�|�d�c�E�0���2��K����)�����,7D����N<X��ĪG#����HӺ.�[��r���nZ�1tW*#��xUq"�)���&����x*�%d�Q�?�%��\��df�!�.�%�Dr5�(�;|�;H��4��"�	 \3|�Y�1Nz�f
��WD��*ypI�:�9���K�:+�W-[6����\���bJtx�R���5�;�l7���Q�YQ�-�4���*[�
;[ks4�a��c\��b:��űE�K>��LS@"�s$��#������UK�xh%��]k�	[�h�e2�߃da�v"����4h�]�1��i��Dhg��=�׏	n4�P�Fs���,��C�@:#փx+�V�&/����*eNF��ZCɘ�v+�)s�]�]ߜ��(��A���k������y�y7�.c=����\�P��u�Ӑ��%���$��x�����b�ϼ�cR�Q���(�u�]�b�9�E?g����*ǵDy��C=
����ż�x�AQ�~S�y�	�iQm��a���_�ԏT{+>�#�|�!��� n_�w���w��ΏЬ1��`�������	"�r�Lz /@FV	�� �O�QԱ�!�ފ@u����#ӿ�rS�e����⿇�C��(|0jz^���餫D�8��nP�)�}�\�1�8���l���s6G�R;{@˰�с(ԇ�7|f�4��=�Sꁝ���s�����G���0�0�XcV�*`�E���Ҙ�~/�;�n�ɋ�lD����Y��{39��[1`��d�8pr� d���C���'�����YQ��|���t~��>!���%{S^$u�
�ܮ���rY>^
������-�#i+9s.��I?/��#���/v�2
�d- �d3Y�y
J+��%NYE���w8��u�L�B�¸#-1�f/���<'�I~!Πb9�G� =��S5�3��t��P�(�V�r��^� ��#˥@�,D���	� :xkv�E�E��<�*�~ڿ �x��=�]o4��1�k����
D,���^�^��y��w�Y�j
cTTz���_��߁rp_@��=�[u�\�eطY���-�D8x�x	:��+f�0��� 6�βS� ��i%q��R���֖{�?��}�ǆ����m�=��Ɲ؆.c�t�Y��7Jj�:��&{��	=GwiF�0_��Ɩ��4"��xXԙ�L����{�S(-���UN�Y׀�ᠠ>�w��baaB��D�&�T�O[�ۑ�����?�H��苆��9�˖I 9,QAg;[��Gm�9(m�N��U�;���^�|Q����An�{��"�T��p��E��*�X	Z�-���WXo�8�K���D|ǳ���:��4҄��;�E���;��(�c��:j²��@1�Ÿ�}P�;�J�bC�+� �7u7-��Ȍ*輥�����Ó
̇6Ϯ8�%�;)���"Gra�6?��!@1� ���."������$�\�����^S�[��@z�R�A�;���3���/q_�u�� `��N&�5ա���-!U�Cّū�zπ��lc�8�ꀹZH����x-M�Ƙ��9Ύ�b��=�.hqe|����8�	f�������Q��:��0��H6b0�'�VHv�%�J!k�Z���;Ĺ�9pH������Yc���X%��*4�a�YlhP�Y���>N^%���&u �M�i�S���!է�6��z?*(EiC�;��0�k�m�-/vF�p �((���&w�[��2�P���'�<��1���B� �����ӵ���Ɗ���)��,�Lk�\�������r��Nɡ���I��q�HQ"� ྍ�M�$�цO�k��s��}��R�B#W�|�7���g=nݗ�~�p��|���
�;aI[5�fI�J6՗�r��dY��7�����GʬE�X[
5e��������Ui��R� ���.�_�����[ ���Ց!H��0ځ��q�Ԕ��Y+R�HG1�)��x�pKB�29�D��q��b��Pr�{S���W��fl^�J�Ǔ��n�(�������`��g�*��/�`#�7�_���S�r	
��5dA�Y��zM�݈k0�r/���&�:��M�O�u�҂,�(�u�PS-�ih�#<��%���dO��ߋ/�w�8}$����[�I�����=����pd�ς�Sn,E"����xyՊ�M\�u!�-�5������i���"���,\AѪgA��0�ѫ��9A.�{�?� ��q�c�|�>���=�/<a�}�+TK�:��XCd���i[f���	�Kt��TB?j��NIй"�����G��3�£��K:c}�m`(QJ��_��2W�_�<��������I��hl��x��D?�%���Qg!�B QnQ{������Ye��&	k�!�2���\2�2���I��)���G��p
1�	yF�{w�oK�G+@(JT��J%�(��!ze1_S�.�a8��x	�:�9��l�� y�t�=�ܵ������������FҠ�r��j���`�� 7���W9J�N�Z���"�Xވ߷mJw$�@>HWž���*�*~nf���(����g�m $�������C�Rg�/O�z&cn�����s�]H�:��ݟO�ju�=����*nzQQ�`��f�y3ϔ9@�`��C����2'-A��OM����� <+�π�W����FԲ xח,2��G���Ƃ���L�������H"6��BRE�1�v�t�z}Ǒh�S�����Y������g�9B��¹�i59j	�6r�xtvD�؟����194U��#��	������8���m���J�3(�Ag����M&�s/���3+ٺ�,^F�z�܏h� v56d�a�1�������gGF�>K?�(�pd������9m�V?�({阪�33��U�6q(-�n�r���T���P"��4п3�lD�KII(M�s��D�H������|���&�7���Wn蟣B�w����.��
�D�k�w��x&��Y����V�8SXa;�, ��X��{:o��<���/ {.��;�}-t����\��j�=j���*b2�"F�n�.����I�4d����W��T��ȩ��� �yBq?#�J%���P'!�����j|\�Zނ�M�|@�T�3 Q����9��=���P�/����-V��m$�Y�?x��h���z��i-ѱ���~f��`A_�@�vd��w�׋b;���+bi��eqOM���I��M#����eJ/*�Lk���s[��}SҬ�~3�I��
DӘ��]�����6$�&тX�`���t�G&,��i�FF�pU�ʥ�ԣ�P�H��yT0�)dV.���7���u�7�YM�^C�Т��j�3��ZZ
�AV��_�5Ѿ��g>M������ȸ�	q{��;�U�	�¡yi���B,������d�K�ܑ�������A�8��@Wu���0�493��ޫ��>��d�&nY�{��Z��z����֤}��O�v�r��^j������Ym��]�������n�K�L������g��bN�X���;(��V+{H?6K1.1��_^���p��b��R)���0�,�߶#'DU�0�p'Q���`Vz~&͏HI�)Nbfc=(�J�=%�/r���"���#�`���'8����ȉ\�P߻R)7��{P׃��2]�~}����������W�k�
�J�Z���7/# @��s����T󾌨��~�x�A҂�5��(K�0P�i��6�D������+ݵIU��݂���`����R�����۴�Fy�̅R[0���(i(m^�����m�bs/IEp�{�A�"�$4�~R��D*t�K�5ғ�'V�)�+'r}�@q3�3�K�RX�D�J�o��O�HfC�W�Zj1�;WT�g�瓒�-b4E��%mi���,��j��)P'�!��"��֪A�ξ�?KЬ;c.�^ �-�>��W5Ǆ�۶��Mer�<B�/�޺�:r�{�K�<�l�6ѝ2��~xB�׻�:�1/c㠓N�����<;�������6��Qp�=���'k�@���sq��9���I0������*#�U���^iX�H���7�m���o�Vb�YN7��O7x����ho+�°�O�FfLF��;���]����b����_Ht����= Y"œ�C����,]>�om����9(�@�|��XoN�ϋ�@��U����fb��1�!���l*�Pl�%�����ͩ���:d��8"C�Ý�Ia>�-������F1z�'7�=މ�"(X�h�K,q���a*�#3��[Of+��B��E�����Z�+�p��,|˾#��%��u�����B͚�"f�+|.��eW.,�?pQT�L�����mO0���%�2�j�]v�� �z�}��a; ���_�/ц|�=,#VG����#���"�&�c���B�F�{�v\Zn��y�f�q6��W+:-}�c�B�ߌ9���s����&h��]�$�Q�,�d��c\����hYPH���7�iO�����R]����Ɂ*ְT
��ɑ��@�[V��Sp�w؎� �ju�u�8�1:�t-���CE7B��6�8E�$���Xg�DTQ���u�슷I ܧ��Hqd�d�$�:�}Аڔ &E�+�b]�*�b�#��_�6b(��vEx�I�J� ���B�P��*B�?~��в�=�����
0O���U����˚��ϯC��Ya~�W��3d�1@�v�;�th�&����l6�pbd���֩E[��Xģ��A*Ţ��n�uy�"B�,�le.�Lj� H8�Erz�Y�D�f�4�E�����<|��]�����A����|X!8ßz�-?�_8L��Z$����y�	�8�����lZD�J8�x��>9�?��퓴҆��`�G���4�>+��o���_sP�I���;l�yU�C+�fdu�7_�~������[%�
,R�)ب6�@YJ��x!����{+TZq�/�2��^zR�(����T��I��L�bSmvWn�e�yz���d(�6Α�A�j� 7aGžܕ+\kx�"��]5�����2�qB."q�?{9󋂅ԚaA/A-�M���8U�[�Z��|��.a�V��9y��Q
лb ��@s��ܗs�t �J�����_j�q��mV�Ȕ�(t����"jA߆�n��g�z?|ä�2Q	�\�ߐ���{<`t�eBʁ$I���c���-R��8���uʺAoq?�J�<08)�J���e�D@�)�ɬ=�y�� Ԉ{U�9h����̦? �x�.�t��FC��i~����Sm���L��y��P�Y�[���J��q��B�v1,R	�E�2ԭ��j8]/	�����p��(���#��d׫h1y�-r�BLFM3�/��c���w�ռ�����4��Yu�j�����'8�T>Pq��Eyǒ�Y/���ȫ���>п)���Ϩ���Cٿ�M_��Y�b��ꌔ,V,�3��غ�Ǒ]�7��+�x8n������z�	䕊<�ߚ}��v %�v�4��#��C<'�aW����Y�ܭǥ�c%Te�޶�ϛ�flV����i�~5AF���s�_�P��@�7T)L��f]f�G����3�w4��t�=t^�Y�|$	K��U"��`#0�q��@�	�l��g&뷴�N��f�W�Xz�뭗2�	�V�u�VX�B�'b�"�P�����\g�����C�A ���8�)M`�2T�U^(B�����lE ��%i0�0'�*��I�3�V��)��5��~q��h��=��G���d��6վY�JC�7+F���#���4-�Cձ}����_b
��|���Y�m8�ye|�q���~��ل�J��n��_X��7��KVn�����=�t7D�:��5���km��O�������)�Y�����a9[024e��	�}�Ʉ`_F+�G鞆�B8�@�.Ŭ��y��ĎT�2��Z%����N��B*z��i6B4��A�FY���l�˟��T?'�otD$�XWOV�9�K���~jodba����k��gl�z]^Z����<�t����I�g| jғ������R����X�[����Xt1}&E��n�� .�N�o7�7
�=*���C�[�|�#���-6�ΖS��Uz�Ki�N^�)�Ӝ�&�lowĶl�B\c&�Y{���\��p"a���U�#/���嫺��@��Ֆ�R���fza��#�xkVU{o�L�0�G M�{�f��y�,�W���w��t�*`U��&���|�AD��p%�M�.�Zzp��=UvǷg�OA�D󵊒�Ң��JӾ6����T��
,(�%i4u�
�K�S�`a�}% D���.��x�N�$��}�e��8��o�C�G�S�a+�"j�#�m��F1��W��k��l�̹��ްVLКQ<��A���w�v�9n��#n��V{3�����%zDC�����W�����"�|�.;�&{r�~�PJyiW*?YF�T��<�L���˕: ���n�D巻Y�Ŧ�������#?��>�I1Z���xT��ǆ��a�A\,a"Tţ�q�B��"�K��La����8�_~7�����aE�����~ds�֤�¤jq0;��@(z���TN��%kv_�����ɗ:��ş��3��$n�Cw���f��W��]�'�%T�2V�qu"�j����X=|b�t�>�͖����9�v���t�i���cط�ҿR��ѝ93�kY��zX�y-	D<$�
�5Y6#㚙�GJMM�;�o�!�a�梁z��՝))��Y���k�XD��Z���@U��h˿��7�R��4�Y9I�U5B��{�r�m�֡�n�{d�y���RV��wmˬ��ճ"�޾e��ހE�23?���ա����
��L;� [���ht�Y�C� �ѫ%/{���Jl�Ok�6l�|s]y�VmŪ�U��Q��R�<
�RЪkr\"̪�7��Q���_��,�$_�δ�*�, ́�G��Σ������vr�J�;��ے���"�t<6��z�,�͉��|�ܖF8��kj��V�lKj�+��:Uy2692al'��ݎ�#3��v��X\hgB��D?�X��Y��0�$��v��g������[��/5C��i�S����u3�� h��:�b������tGE��,<��	[�lBЀ�\��ߗѝ��^�cc�C 2�O!��h��e}�͓�ST��sl;�� 1N^�EGT3|� j��a{[SVh�OP'I0�[�`{�DȰ�p�_�v�r��̎�)��2}Þ�ba#yt�B��N����0�JFK:v�|N$�6��?}R顎Ύ*�����0�qh�� ��%�!��K�̲��,���	o��͒�����%�6#q��/gN���/�
� �mm>..m�7vP�q��&^ǚ5��`���qL�\n�qD�DS4��ӵ'݉�19ꔢ��H�.��h�����[\)�d?��%���0Pe�ܷ<�.�)G�]����j [7�͗�91~��1�щc7�it�bյ ���3�vi��td/�K�����%� ����s! &2:sA����`��y���`Zh���3 ��AJK�{�b��7��TpL��t#���=W>��F��޺R��l 6HZ]�^q����U�	t#�e;x9��(_��|=Sl,�b�ŸM���|��(����zy�k{�LmU�r��0�0�7ȯ�u����q!�}�F��28����!)��%2�S�V⌲f#Ɉh�H�������G���B���3%���sG��tdX���|��>C���p���nwc��u�>����H��5'��?�M�W���NZ��u���{(�t��$	1�M$��|ߋ�������n�"ﹴ.ޘR���!m����&������}gQ G&фV��j�� e�� #msZ<��M�K�ٯ^vק�t��]8�7Dl����m��ݫ�!7ȶ
��Z��� ��a�����KA>���}U]	� �D�/�\�+/d ��*G�R���
���P!r��:0��}ρߡ$�x�0�t@-��[�Ʈ�,>�r �!�L��!��4��aRٶ��i*������5��c���A�u6�v�M�h@v��&p�[�j�������I����g=��V��p�N!O�B��Q�V��Q�A-W	�Ij��dq�\�hf��;{���ӕfvG�g����<�Te�-�ӧ�)��#g�3Ⱦ_�'@誦�܉���,+\����e �������,�C����̎�C���х���3�� �m�Y��f��s��H^:o���Ug�<����������h(�u�"e�Uz|nF�����Jv�Fi�	��i��W4'�x@���ܜ`%���(�]�ػ~�m1�y�2 ��]4df�),��=cu�:0e6p����i[9�괢�`d�����9(�]p �;{�'��[�^Ӯ�9��?b��	�����=����(2���CB!�Т�3i�*cV�9������L������XQ��b��%�x!�t�'���E�t�Er?�n���*xT�z�ҋ	R�`��t�=���+��U�~���}��7/���0�f�^�8ln�(7�KNP$��Żh�n̯���n���qv��f�1ګM��|�6�� n��Hdf�i<�O�[S�����X��]:��Wt�s7�߰��ry��&ݞ�X ��}��e]����]�A�q���!w}�z��
���Z8���L^��.��SqZ����m�~���G��ٹ=�'�7���������7�#o�c��B��h�8{���ա�=�.ֲ&�ʀ)u�h$�Á:�/�"%�c���-H�]��ݤX�n����<�Mm�o�̈�2�RY�3��&�o�ʲ�L���I*��#+�$��ް4^�^lӳ>3F3'�.�O���>�,������X���	���iTZ(=��dսx'g�9��)Ѭ���	"�7w��5������\�*�f��ڣo�=P�A�6V��R��Nz}h�(���e����S)]>�J9x*����a}��VʔD���~��R9���j�W����~��I|]&���$���v�ޟ��^ ����B�g�ķ�z�l�+G8|��$v�
��ǻϢ�P-(�_��H�M�8:�[p�K�%�E���i�ZG=<c[�9",����dY^�9��|)i) �d�\��L�+��A`��T�Gy�F��An�j|F�x�#K������[��Ϳ,=��Y�}�'��ƴU��@R��J������-oM�,z�'^황��z�Ւ���F<�e����y<�]B>T����@,I��GWk1�7��v��%�:��0�����Σ��I�n$�F�%idb�n��E��� u뾞���v��'z2a�`d���gv0}��Sy�q%�k�v����b����a�7[	��MG�����o�'���nr	���-~
�N����"j�6lC$�|rؾ�%#p�ra��3�(blz/���=���P� �2��"��+���YԬ���LM��)��`GF�9�̀ɜ�y|5���[e�� :�sf�l�M�R-=�y,Jz���m^�63�v|�q&��=9xv�L�ܓ�U2���Lȵ�R]C���ҩ��F�%�j��:$�r�}�)�D�v��a�.�uev��8�I���'>
�[S��&sIp�g���1�8��/"���	���C㌞�]ٱ- �D��d4�ӟ˞8A����*A�� ��il��ҊHｺ��͐H�pY�.F�G\@K������>qK��U~ r�=�����R񰲝{� �uʢ��(�#��.]m�4��&�E�� 1r��Ǖ��}aNq�e֨-�Te�@O���j^(���Æi��mt���l�X���A7�~+�8[?/��ʈM�<�=�s-�3�*�A��3�	�O�~�C�K͡;y� �l�(l��G�����0�n$��8�/D����:�k�#	�o5`@���P����-�=§��F��z��h��6��Gq
ߗ�f&~��|L#��1�$�,t��C�?c
���c��%�����e���t-'��f��7�8x��}�B�*��	�ศ�p~`Z?�iI���u2~���쥑�w��n����ˡ"_�oK���䕳�����؋S�r=\q�z6�R��B�u����8�d�+���&>�U�ڨ�
�p��n�qV�B�R�L;�e�?>]�r���<<J�:S㍃��D�R ��xd]#<sa?(��S���p�^�BD���l1iD�L\y@jQ�����/�$��% $�4&|�_��2�Cuq��1��+j���=AX��jZ���FY�=GE��!\�zD��@��C�z9^��#Ð�٠�~ p�j���=f\�I�:�����6k�<�T�����<6̈�N�	�Y�
5�~��}8g.g�nrG$����/�#y"�K�IOs��a��ɷ >�����M���;LtWŔ�M$H^u�{b�_����i��aU��O~�i%�<�0�c��0(��eK�,�����juk�|ǧ��Cl�b�bl;Oe��?�{\�jˑ՟��s��r �I;-�O�d�l�	�e�l��!fח����mƔ"o`�y^_(`�cƀ>�୭��kWh�Q�}8����e��[-��µZ���v���#�2�c��0����� +/;*{R��}��%�g���g�o<V�됫��>����Y)-%����Yv�]�2hӧ�ͯ���u��*,wN�}����<[`#�����M����y���i;ŏ�ȶp�
luBc�6ݛr�K��(Ɛ<�8���kl����8u�&Tp��*���O��W=�|���h���mF�*=e��אN;�Ҋ�T	��b��[�<���g�v����`7m_`#^���]�
�rT�h"���;ϣ���( �sj��Gv��Hp^#ќ����U����k<Zˁ6W�_ʋ���� E��"��O�(2�LN5=��3>�4���t%4S�Ld㟄�����x�K��[�r�S��Q�»W?�KB�\\���������X����x�Id)�#x�7�}QȬ��d��	W������=c@B�0�(!�j]#e��$O�_@cZ��g��K}��7)��@�����s����Y������9|� ��0q(�E!��}ן6���h��N���`��`���U���f����t��.��GZ؆wr�j�)@<�t����Apg`n�-س�j~t��]ƜN�/��0��YB�96��]�j"<J�^��q��)���5�]U������V/[���m'M�%e�N�-�?�y`�'��K{��s%�.��9Mi�G��^�w�4��K`n����0�p�<��7�f� ��+U�����O�%��E�!n����V�/h$�������2�= ���p˅+$z1�v��K�䌯*��+(���6��A.E��4f����F�4`I�:�hM~/Gk�>�r-������a��]����b[@���,����
0^T���1�^O�C�%��O0�,�|����Kd4_�>¬4���
R�LG{ڹ�@<iң]$=�c��������I�h8�P��C����ܭ�nY����.��5>�q5���<���J�Q��(.#Ȁx�òO�����1'0�?q�W�_d�݀�%M7�ז�����VS�z�63J3�k����=��(���*�	��-�W�]�U��`�Ո��p����?&�0�j�X%�H�{9M:���Lk�p�3���Cҥ-�CDC��-��P�R����$_��u�lC�pJ�uFXZ������&��و���dV++8���)Ϗ����WP�\c�O�cN��ӽ:���벴�������h&3���� �!dmS g�`����/ĭwUGr�'�;���� �Z���Y�7���(��.WgC�t�0�`쒳ݨ�TL���G��p$���2�ast˽���_�(����U���B��y}�}�_��a%���f=��EJp�Aġ<�ڮP��z;��~�NA��u�b����Ϩ�T�2��T�Kn��&�I�%��TL�`)���/�<kH�� Z�R�2b�ZlB^�K#{zua[]��M��@۞ƨw���%_��R�>n"�b�>�¥?cT�ª=��O��yI�3�1$ar+��4�A�&^"�7���}\jW)�8ޏ��"��wo� ;��U�<���H1�ޟ���P'��b-g��Ľ<���hk�:�[��~�<:��1��uA|�/�!q)���5;	�p�	�/�V�1u!�]�2��R ,\���F����'�@��U��*��%
�M<^���W8��~屋��)I~>O�{��6�b�xB������U
j���}u�C���5㵨t<�4��E>�9�l�<���-+~o���NT�0�3��%o��s�AK��B���߲?����D�k��PU`^�
H�?�z�������88�@��{�l<�{�F�|5	1ĸ4e����͛��/�MG����r��Rᑏ��ҥ��ob��U�d��B3�o4�;��	B��d<��E�)���9{w>T'e��������L7��q]G)�5a8U�n�>>����D�u��x�ms���ߩ�I��]��!�tv�k:j���>h��"�����k!j�E}�o�(����'��O��4�M���ͮ��U�s�±�~��k����9������^b�hA�h.�y�mm���#˅�'��f�:n��J� ����5W�Dـv}��45�(���>��J5#� ��g���WfT�E����oq��t};Đ�$�ׅ�`1�3�m�9'��+���>���0�H� ��{�r�����.� � �$�{�����r%cַ��7�P>��F��=��H��A�dG���g$�����z7�cl�݁E̳�`92R)S�>�.e�#�o�g�"*:M�-T�Z�_�P-H`�1��W�ɚ"�hg�\�����"|��5n�/�<������&�qz5�CXL"�(�y�p���JRξ�%yk���]���:��'�d��*���X��7��k |�g�������@��өq��
�b���H�\��I�@NdI_���c���kuP�u�Z��F��si���r���u���>3�&� _$}Ӏ�F�a!��1t��A��p� -��ݸ[}ޜ�{.Ԍ���KD�'ي#���2%�4}
[s�iY�����q��Y<?K/��k����~]��ȦcBxCroO�C�1%�ס�z����-n��]3����b� ��T���9��U�
�*��ι����5��8|������VY������C]J)Jk
p�������<5(�v"�̒?�^�O����PN�E7:_���W,a�P�_H@�5#��k��R
��=� n�46wN��~c�+Kb��܌}��9�$�������±pz�~)j7��,[��U�	VS T��y�K�ϩZJ\[
�B*Ē9�iZU�c׳R\y���X�?��9@ߺ��!�w`迹��"�A>��LG;�]�D�c@zD��D ��5j��`�KG6��9���#����%a���E(�^=̝�wa��t������{����Q-���6�Z�-���!h� �̕�n$�Z�5�w$e��T��#H�����1Zh`fJr�N1A�m����w_��_�hȮ��{w�F�&�U3���ﹲ`�氊��\�H�Y�#�.�"���������U�"h�3��`8R �=�'����"��Z:I�Ȃ��R��X� ���`�_t>��:2���"�
y��̡��>&�ћ������{�J�G��]�N�R������ӡ��{�"Q���V7ɜ~�Ns�� �c�~��Vn��C��"�0���2���2.F�ˢ��,b2�!�T#�*� ���S$��N��]��ȤƗ�B�i�F����'��"�V�c���]Y�ă��|���m�aȁ'Fٵ��3F����
a-v�����W���S7{�lp���\��#,��Go����ҶUs���G���r����~�wQh�X����I�sG���ɻH/.�u��e���3Ȧϛȏ�e�����i�ikW�� �$1�j�~��K��~G�$����(_Q�;���#�ڽ@����,t��=U��M$Wq�&'��Y5���"�u@>��0���wE�˿�s8���Z:�:� �a�ߣl/n�f�ZZ�>����~��~)�n#�>����L�;��)�됯T/�5ː��3��MTu&���~vnD�]g�>[6�m �+4�sp�Z�i�T��ǛMϳd�1o�_g��Yȗ���h�3&���X�� ��Vy��:νcvBf���d}q~7����g�KA�=%�ی�4tt7K��@�wT� �#nn�ip�����&R�'��6y�ځJ��ϮP��A��sR"�g�rI�ab&��(�
�����4;��L%.�����O�� d3}��N�JE_���"7LI�?9
���*�D�[�c�[|w��R��
[���M}�s<�1�A����0�u���t��߳O�_;k��mΆ&�߭��(PR%�쓽Q�+��R� 4�i�i�DiD-h4��7����N��=�o� �-,'���v��1���|!)�*:$8���?5(��B*O�����x��b�h������Um��1��d��m_��\)������Sqǔ�`� AwA��HD@�[�y����ǉL��n�4�I^ �Zr �����/���y�e�=��M��_0��[@��D��4?�k���(~긺ؗ �oW��x����yN�&���:9|q{�����	�+��}��c{Y��a��?�m�}y�&�X�T̗v{�9'oс�x�
n2�Y����8��VW0Ѳ��j��C	�r[�>h���rT�N��W�N��:��雲��JqE8�1��ǸRO� �3��������[Y
D[�e�L�\��Kѐ2� �Ci���آ���Fbj����Z`Vo�,�1�9;�
���ڃ
32�N)j���ٻ�z������'�7uטA��o�j��J�K!���͌m��o3ߓA}pN~�N�'���
�{[����<���+sc��h+���^tƚJ��s��~7�����F���Yk��f�A�T������m�v�,觽��[�ً�FƁ�������^n|`�֩�W��DJuKgFt�y�|ܻHJc�h��}�ҥͥqN�;2K����b�oI��0��Λ5&3+���k$l���C%��H<1w�u,'�ϖ��~�����<'f	/e��(��t	'�r0�p�"P}"��9�|��{yk7�L�i��S����	�%$JJE1�����4*�L<���7�Q`��F$F`Ǩ*�<�2��C�u�W��m{�h��}�����?�رٷ��8I��� ѿ��"
^����g���'��6�hHpt��?��_,����C8�, �4
~꽓\r����d��f[]��U�qk��Em;$�U��A1��Vk&�~&9��O��O�Z{��Z����?��W�n������j�j���N�ĸ�A��I����6����N��|�#�{逭hˮ���1.R���)�	��f���j�x����cڥ�k��ڏ\
��i;ZS�Bd� ]Y����5�"߇�� �x�帥�� ���?���ڶ��u#����G+'��2y�aZ�]bh#N�`4�N%/���q��N���_g!�X9o��΅�8�Sg,�k(�Tu�~�<���9�������ŽOE��J6@��t_q:������cɐ�6J܃L?�bN���Y��?C��?�֧B`�F(�&�U
hF�Y�0�daU��%�rW�����t�]�E^XĐL�z���)�.:k�=�1���j������[����4��U�^��ծ��*y�.��[�VV+t��l�O��O5�>z������ٟy`�T�i�Io�9��.�o
<@�ח��ߣ��!��B�9IH,����x�\Q�q]/o�Í^[F�G�Q=�I�Z6�P���2 =���Q��Dm��.a����6�/(�4j�+C�����4~Խ�ՙ�R�;�܅S�d�MS5�6a�]o�dC�RԵ���{ͷ���_��Z�=���y�I� iX(+�L�.^J\0EK��~��fic�h���C؂s�7E��m�}6(� 1���b��|���k�}�}�+4w��՛w_�
����+&&�:��O\ۛ�6�Ѵ$G���/����I&}Go�HV]�z�ı�1�.h��d���ZcZS(��a�����E��Zз	"@�H*��.@Sj�+�ygn�މ\ڤ+��v�>�b�L/h��[���j�C�\� �O�\0��A�ah�ZZt�	ec�0j1�_qQ�	̘];e�������P�\I�����6�Ǽ83�{�%ޫx�������'I驗ec�,]Я���?^���S��7�H7�����7��1RyW�>�K������e���]�e	l|�����B�v�@���!�<�q4�+�Ļ�ud������)B(�k��/�RQ�c���X��!5�ɠ�|D��W��vp���G��=D-Xǂ��K�oZ����&���\o��s�.�|�wam�UL��&).Gs�;���+.)�q�e�U���	)�F{�w�Ùr�ѹ)�[�ٍ�4�tk̫�{3��]�N+��t�����捦ɯUu^}�\4)��"�Ʀ,�+4�n`YT�����m�S�&�l�f��]�u��w7�G*<��ܽ)aL2E�^��41�mo�ʵY�w-��<A�P?�a]s�A�3��߿��%�b�t��Q����x*n���� 9��O�3տ;\Ίyo@�V���b-퓼�G�ɭ$r"�A����Ц�Q���B*�!���R�W<�W�<R$k����cGs��A� f��)���MX<��Z/��;u5T�F ���cf�߈;�u0�*�pB�=�tʚ@���}5�N�"-F�LZ�X�3,xv9{T� 	�ъu�r���T0��h�t���s�o�]�V��I"��5�4I�V��;�y�C�Q>!Ņ�շ<ɜR��/��;>���,Ș����BF�nˑB������Q>���3c9���`4oPu�|&�H����;�m����F�D��׵�����b���������@��*��֝x��"GA�;��%��E�����pPA�V�(�6"��Y��?f���z����k�|��0S-W��N�x�ݟ����g�_:����?��y��Oʵ�`Cu��C��3��6�o�$��[�z:�H�������2X��jU������ƪ_˂�����?9S�
v	D��	L�ϫv���oNQi��Ҫ��>�>���w��Ui���VOM*R$Ԕ���3��Z.��b��.YѠ�OM���l�F����"�9��@?�N��A<LqV�����2�Z�Mm�<?���U��L�C��K����	�|HyęS�(�ibCI˷�*�i��׾Y����=��<�и�Rx+�q�v����>]Z����]��ڜL��IP��x�[l;�FBl��ęO�p������Z���L;��Ή�2���J�jb�XM[��%��P&��M� �@�f_�m�FL�U��n2 <�c�LX��j7�B��y���7)���)���Kn���%�����c��Tl�%}?� ڭ�(�EI�qۺ�v	�
���@��Y��-IG�f�R�,X��	�ƹ��C 73p���0'�����f�##
�I����zR=�_i��z{�4��+,�F�<i��N���m���]ѣni�=����(����RJ�ݪ���ILo�6=YA��ЗZؑ}K���9�9f�Fe)D/�&8���>l�"�U&B^�M���h���tZN���*``���d���/�S�m�����0�OL�#�r�:,�*�3t4N
E�]��[��gD���!���ϵ.$ؑM��������h~A^��s��v'���˙4g�uf&�|8cZ�iw��H� ǵ؁㪞�ɉ�B� P#hx8-����܋�s
�S`p_�l�.d�����4Ҕl���8�FK=]`_���XT�I���^�:��:��|e�_����(Kk�E����[�|
���n�k �2�Vm���x{C�J*D�Trq�� h0�K|�ƺ���y]���V*H��S����jN��#e���=��IS��'�#�v��Z�4/D����k�B ���ί!�t���=���B��M���jD�,e�;~q ������&�)�d���ig�c���݇v�c��tL�\J���<�ʿX����A�=L���nr��V��ڍ�����΀�`6�V�'�E��߅m��l[�E�k�_V+�/}�~%�=n=�%/��`��[�w�!�� Q�W~�(�ݧ=k�u�q<U7{�\u�	�4�{��؇��f�z��+�wɮ);=Y��v���ß</8�L�*�&|�wF�+����<F�-%�#<o�I��IC~����
���,~��H}��]�����(�l�x)�{�²�B�z"Êx^�����c�AM��X��k�x1���`<M/ޤ�p����_��A���mE��]O#7�s{!6��C��"�a�ϕ��fK���}U���om�O��Xײ�ϯtf���M��a4ST�7B���H�'�g��y̗<�d����c+å'+��c��Mh�M�=Zͤj���-�ۨ��.�&{�I�ǽ?S��C �i�8oQN3)aUcnVE@�8�rM������3��/�� �ji��.͚�"C�Ӭ:��2*��AV< ��u��4 �#$v�B/уA�B:����<��M��߂�˦[�7q4"��_�p]3��v�*?�<B��qw�B>�'�@�̚��e�Q0-xM����:�;���Y�'�A��M���к�SҚ�ʻ���:)2���DNw8��&O'[/�=N�ӛs8W�n��4�vԈp7:�5q��h�#��T<^�8�Η�I����ύW/ǒ��zW�:�kw�`.����zp�"�Q��!��������Yz��8��#�a��"Aǔ���ۛh,�
�pu�%�fC��ߡ��%L�:��gY,U�w!R}8���ܝ�m�o�;���(p�A�Q������s��
Ln#��`蠓&eX��]k"=�G=I�!�4P�v����_�F�`�.�y���t��"-�va&��2�5�4�׹��3g� �&D�f�$M�c���i��c�����G���{w|y�[!�xo��T9!��D�'6Lܵ.��M�\�TU��t��T���[�aM��z0,��a�eo�ݕ�2�t���li�D7�<N�_-�5���Xxf��&��aL>�aEK��S}�јl��(r����e
��K�\�knu����i�/�n98��=���½����R*�H}I������|�#U��w ��}�Țg��`��	�rZU:U�������څ%�g���T�j�9(m��L3�]~c�&�I������,��=6|�J�Fԯ���d=r0�.��������v���`��>���I���9@�+�
�T��#Yx����	��1uRb�Hj���n_t��w!�n�� �S��¶��eL��(bUu��Z�}_sK�sr�y9l4^鴂��N�$ ��M.��*�����ʥ�)y~'�%�����&G����?[6�ҁ�3}!�~��?y�=P'ׄU�h��:q6��2�?r�SR
�d.�|���Ĕ2�_ޡ縻(�h��Q��m�/C��֔���eb�W2�""_;ZR����N�^<`�������6�R�����l	�� �w��R��
;(��y9�o�~n#񁞀 >��р.�j-������}Jd.ARylvV������o78XO�k�Y�N����7�!��U|>�j`i�hj:'�?�e��F�#7߶������B,?s������m�TnRP�ӧPC�\����d����N��mjų`¡L�+Bz� d�!j�:�^])�w�K���?��֛N��ڷZu���e~�+���`P�B�{���<���c�x���N(S��u�{�|�W�� �"?7�Z��7�u=]L�|-��dB�ϛ�j{�/T̉8�B3�V�oQ��I�֌�L�����ֿ�(�
���K��,��^'ǥ��m����q��S�6���CV�����e�s\����dCa�w����������h;��X$ٙ��07���AK
�H��}݀%ij^�<Yq6��B����վ$���N��wz�t���ň��ǘ�ڧ`F���Z�l�j��~T~�'0�p?��vL��0d!{/�IA���m����m�W[BW
h��S=@WQM��\�����ч�Ė�y�R�`%đ�|�Ԥ>j%��0��x��AV?��ϬVɲ��s�g8�q����-(�Ꝧ����G'�!�ʓ'9c������������1A�+M�Q_�<t[������<�|��wa5������D�8u×^��
�L1���3~�3�1�X��X]u5�������>�e���Fΐ��7�Wi��U�eE�g^zF�iM�D�w&ן/�w�vɉ���X}o���?�X��[(���6G ��:I2)PEoF90>)Zz�����"Twث��ĉX�� ���-�yd��Nu�]������h_�$�lcB�@�c�����i%x�I �s���V�Y=X0J��A:�"i�iנR��a>�w�1����_|F�����zo�*5�����z���$��/����|�tk)|�o�A�}q΋B��.R����5�����i_C�S(u?�WO�cF�="C�3��GEd	��(e�Y�����#��$���7@H��ǐ���SL�qa�;��8R�&ճ��rF��U?���;� V���WZ	�u�ŕݶ.�kL��o����Mm
���J�g.���K8��:,+�T�����#��F����@3g�\`G�e88]az��YR�r@��GW��Lȟҿz%m��p������z�#�E��!fv[�f��}}95F�9�j&��%��E�&嫧��͏'���Vq��_��`�ݡ�n���^�}�A]1��r��>�H���/'�K����q޹�׭M
.ޅ7�SǇ�P�A�4���*��5'�M	�v��2��C�J��e 6K/�f`d���xw[�L7�Ԙ�D����:/j9���A;�݌�ov����=�6��c1B��~�I�ˬ�ؖk�g�"ߛ�(+w���n�n�ݬj1��שs!ǔ�ڬ��&N��Q�������{��d50mH}ms�
��n�J�)�3R�1��-^_D�HO�o��ʋ���ֽ>r�@K�ʀ�� ^,p�(��+*��	ms��������^�����`��=���}]����HMZ�ڈ]:~��S�U��:��¥5)}��[��,�YԠ���ϧ��l�Yf��4�U��*h���:��4"kv"z���dP
w��m%�Z����Q��!|���h���}����1��AJVB��/n�sbf �p���e�,fC�>9qE}lfp���J��V|c{7�ͪ1�R0e�ƃѺo&����A#�j�ud.t}x�05���@��1`�b�"��L4������mmr6t�8V�٨��.wv$�l��~�y���
V��`m]C�>���8���I���6��Wr<�Ѐ<�u��p=]�Y�ϵ4����J+��^���5�;$Q�߂5��~����0;B�~��3���JB@����)����{�\މ��/�d�lf:��[���ttm/�����g;rhx��[3a�+d�_;��Ф���Rw��.7�3v3G�k+@��+��k�z��u|���}�!o-A��w��S�y��2$J,�ݥ��d��5�]�����4
�|�m&��M/S��e�b^�ar��O��w�¿ф�8��7�-h���	��2�a�=�Ox��3��[�YS ڿ)W�Ş�6�H�83�D�.�M�����X���٣<mQ��0[Jf.�Q�C�|���å.���Xkrhg����qNS���5_�F�����&��f�wI�����xz��K�3;7ƛ�$�e탬o� u�6��m?K�c&e�{�xX6�zh�;_�EV��U-l�l�:ZX��XW�����~4�E͐ɔ���4횞�)�B_lꗡu� ���]��n{P��w�L�
�Q?ݭ'6W��Xo����n�A4$���&n�SC5�b���[W��%1+���e$��
��r����[;Ƈ��PIA� c��3Ň�+v���V�=�"�����x�:����2�	�֎yw7 ��NK3��"M��AxPR�x�;����:E��w�j��=��b�9ՕU�֛g�B�ư�')����lOп ���~���@�7����6����\ƌ24`��
�����-�Ӄ�@P��Q)�I�ܾ1q�6���p���F�޷7�zX�?mޝ�J38�����)-��u	Rv�µ��a�}��N~$�ٺ+G^/�b�*��%��i���׮q����lX(Sm	��9����8Dqڞ�8ߤ�����"��'[u��ǋ?��ҋöo���U?1i�
2�zIH�������T_�J�5���P`��e?��_+�L�ם�F�o`�+�]�Vu&�EXV��A���ŗ�\�A |69�kr#�R���̭�P]T�bYQ��Z������E�9aJ�9d�w,�PE��ߪ�]8;����F�h��s����E�|XWC�f�$]� �,��{���'��əƀ{ )��>
B��$�C@.�Ft�>)v��=l�[FO�c����H�]sF�)��Ib~e��CcĴ�A��66|��jʨ�&!�i�!��ݙ��b�
i[cA���A`�E5�*��	׺�~a�;�4�@?�?�?I>�Wb`M||g.�F�C���[�\�۬��x8�~L����;  dL�E�WV 1�Ϳ�}ߓOI3�r^`vx� ���@SUKat(OdD��W�dQÛ9.9�O��vT���>�,ɉ�k��y��� @F���i]}c��:��lp�;҄��4o�Qݳ��C��Ib@Y���:�c���y�u����=�E�,���vT�M���|'���;p*wt5w �7��ˠ�m�(6q�M[�L��v�}i�m/�mc�l7Ǧ�Fw�^)Z�U�]PO�5���,���5hE®��\A��\��Is�����?��q��zC��+��(��?[;w�����e�C=��&��ջ�Z��,���;�H1g�e �kvɄA�5U7�C|@]�cˉ���?������W.�z�q^�!�%!��x-���яe,MI������I{ �����gcSr^�~zʂ���׮�u��%�;������FM�O}x��.ظ�����)j�+i�f��a������ �Lj1����/a�+|�p �$��R��.S��ƹ��g�4J�b_���>��!����%v�<->t�U�*S&('8����홚��-0�g]�X�j�����aEE���%�5�a9Y7,��Uқ)��^��"O>^֡6�)�6&2�ފ�=z"�N�J���=�����↺b�	���?rpq
>ٕ��(6��=��[>�� ����A%&���.x���	��z��ݸ�2�=�i�c�ȑ���R{JT��.�$�7C�Ȣ`	���2A��	��_�1آO�M�1"����_ht87F�g���IS��a�������mћH�haq��"�M囬��T�����{qUG9�>���N&">'uT�Y�f�vO������ܤV5BT3"y�c��?Qi�7CE�[5�I���G<�뻅�~5�
�l���xϚ��_���p�O�}\��8�>xHXGA$��J��8����H��q;"�N��Ɔϛ�a^�P��T��ڦT\b093�U�^�Sq�ٮl �,�b,�֭�Kx畏! �CZ`��%�1Lh~V��C&���O�;T�Y:�2�d�����]�p�B�5!�?T���&�$����QC�+�Ї}T�F�&�O�/Ҽ�J7B�$����n���Jɷ���Ǖ�5����sA#�Z���O�!��87ny�{�l�����=\=�`m�0!`>6ho����"��W���^!�H�t#��_k�6��s����!J�E$�gk�1lK��lw'(Ӡb�q:�.{�RoI2/{�)��b*�9����)I���Kӻ���d	@B%�Ymgԃ�=�&��������Lo є�A��OU����	���_!-�;�c�˗�0�P���!�Ѣ��@�0�WY��H�i��8����1�-R�n���1IW�2�Z�풔$�}u���П�`�S�6����	{<ߛB�G	r��x
�uq�3a[8�(؟\��[��b�,;N�:*i<�ڳOI��͊�x������!42�55�R8h��1�� ��zU�+���2{���x��*�)��ޑ@���Xf2�U?E�L׮���΍�o��Q��,]!����^Qj� u�6�6�(��a����e{{����s���)6_��U�:s�>uX�����o����K=\� ���HpQ����MB9�h �Q�E">da��X���ɒ��|p��	��ؗa筁3��e�~cU�9��=X�z/W��d��8�f�Q�:`��&\�����#�X���8�ڲ�N~ʣ�����r�M�I��?�}K��V���nc��Y�u�c��ؙp��׳��@\Hg��Iu1���hZ~���a�o�D��ͮ�S����˘�`�;�   ?��v�:f�$�*
\��K�f�����WԌ׵>�4���EĆ�f�K���-ݎ%Kez��T�Y�~����=���S����]G���u���5w9����Aޕeǧ�x�ز%rOL8`(/�#��g�[��uӔ�!� �K\ȗ��μ���|�)sqZ�1N��}�p#����MA;��=_�F��}k��T���i��ޡ]s|5΂���iձ��s:z���rZ��8O�7��6D�8g.��^7��P1)�@�~:w�����Q���Ԧ@я�k�$�1ـH���^�-T�+�5�5G�MUL'"��9*yv���p�;��:a&Ѓ��sl�G�S�V���;6n���Ƶm���Ծ�J�Y�� �*��Ɩr����v$.��L��D���D#c�-���:׈_�����������'滵�w7e��,b��.>h9�$E=R����u�5������h�j�<����� �IN�0f�᭔��(�8U��$�z '�l]�AQ�0J(���H}����%=+o;����]u��0,)}�_���4W��/Y0 ʉ�p�<cߥ�	���UߊrݾS.���G���Y(��1 �H��oE<���^��E:� c��~�Z���kS��UN;f�B�T�2���Oq|%��y��-�b��W'��Ex4��K=�Fm�|�:j(t�/�<:�|�'S��Pb  T�u^?��8�#��)���o;�&X0u�5*�f��m�A�����DP�I�2a89i��QvR�D_��a�.��QiC�ה�_����6u�(�YBW����S��W��%���铸�0�n뼜���ԙ�m�>�\j�CwI���|��,�e%;�_VesJ4�{�X_�u��k�o�1>)�q��}�1�j�c�n�i-�8Ս`t�0Q�G/�0b���.Zz�05�\'NU>=�6���q����xtE�/��I�����
����L�0�5BU�mw��͒Ƌ��`��H��S/e2F� �� �0��6���mK��n������،�����d��-i�+u�'(��J�۞��3`з�wX�� (�/[B�+s ��h-Or���Qx�������$2d6�FgK�G�b!�t�{�$�ek�9L�>����F�E4(&ȅ��vpՒ��
���[��h�����8��(�g6\w?�r��U�g��7O��UnlF���*��(O�q�\�^�����I�s����JzD<'܁��V�Q�AdH�W�	�G�wU��#/�G�,���9��eE�F~:����U�B9G�;윧���M@"����Ђ��s���H� ��c��q�Q[�m
���$���N�"DW)��	qn�Z�M)�9��}�Gsv�_�b��|�Վ<A�5����l	�Mg�޳ı��h�HQg;-ܝ����\�J��@��V�2����x�p���/��1u�QQOBG��'le���5��p!���z,<mq%�	Z��b!�>�?9��7����[����w�ra�������ѓ�y�>��p�?������a�y5W�XM�v�=꤅��Q�����4j�2�qG	΄O�:4�11���0��:�2s���w��4�Ǭ�Ӯ����B\kyd\��_�$a`Jn���=���PO�ؠ��Ԣ��b�{,���^X�Y��մ6�
#'ʇ ��QT��⻙�HQ�^v����m��_� ^���<����ɜ��+�z4~���1Q��R��Z��r����u;����cGSf���Di��1]��}��d�R�"H�ڹd�c�5����X���<�p=Ś�Q�)�\��0�m]�!)�$@�W�F�*�������e�ǡP��X(Ʊ��"�@��J9e�o��ħ�rTت�~�j������v"IV~�a���w>q�;ZB5j�V�鬟�x����n�7	�ߥ��ٓ*�}�͛���A7�����u[D�?dN��/�����Z�{B��Է��i�ے����yc�k�I��~���m��l�.�K�7G�j��I	v
A�j]>��R^)��&P1n��{�tJM5r��*g�l,�
��3���H��m팞l|���׼�ҺxPrؗy��T���/Y������[ 0��ݷd���d��#F�B?zz��ܘ�ʑ }N�73s�M�K.����JV��7�H� ѻ�'[{��q]�|uͥ�d?d�ԫ.�"!�$�Z	؁�P������ �BW��C����U�#ز��x�y|q�v����~�$��O�.Xh#��["�����N�q�t�}nn�A�'�2s��A��8g.���|Kpw���,�R��2���հ�Z��Y��@���M�g�/����Pz]���6����$#�r{�ɉ-��w�e@�}`��ߙs!���O�=;�eW�y��1�A)�,zً˸��%3�͠�L���z5��&��J!�I�	uB��s���,ϝ=�}}p#[ϡF[�.3����Mw|���_�Y�?����7u$��l�8�jt�[e����ACDv��ih��O�h�+N��M������>��Sd-�R�5����O=��ry�r,�Yx�L�)'���`�ѽL�Öl/I`S�]�ك�\钱^Ȏ�Z�ꈹ��F�P��U�!S@=:��_w�:E��L��mv:�;L;Gݙ��+]!�&����Ħ;���4�T)\�{�<}����Q�ڢ��P�	�k��O��@�L_a��>�'=XG���D������.��U���
 ��y�o3�!!�_6���q�I,ތ��� Ͷ)�IhX̹�����iW� -�W߰Y���	?6}�mf�a�g����S�A�%xҷ�"ӈKG�~��Җ��%2T^Jpi����2�%'Gl�O�
.�0ЙNܐ�=��87t^+f�J����f-�z�|ANM^�����ڜ"#�����O�fK����%bk���M}��zن�r1'rW���J
�w+f����zZ�ΥU��O.l�ѭ����v��� zFu�E{˴�W�殽=yF����yq'n't��r&���W}����p@�%*�ĉp����W$���Nq�d��ǴR#�H9V�Qr����Zt}���O�D�y��b�c�Z���<_�?#���N���t�t@�(~S���vT�fʊ��
�TF�O�� V$#LT�&��"+/~��:�j#���K��"-^�m~��!�Y���2��'3�4}펠69ä�I��͏3 ^D��./��TOx�b�!�?�<�>�G��lE�אg0��ץY.Ty�0�@��%@2q�|bGT�2u:x�o��ԫh^{��Q�S�5�|]���$t�~�P+5�ڰP��K�!���ir��[΅��eL��ȓ�Z(�7+S�j{� ����i�M$�Tº������T^$`�S���Ŧ(!f����y���m�W
����%.#�Uq ��Ι�3���s�|>�]N�t�Y<��C�p���q4.�d���s����l��
ہ��q���i������yn�箦D�_�woj�Y���U:{u��1�
�=K�MӇ-�z�_)v`D<�-A��h�@Ё��p�*�3H��љ���ȗ�J�o�m�=����۲$�]��+����m)�N��Q���]��
�<��%�jH�a���*��ǃ�#�2��7�Q*׈���<����+d��Zqk䓞|ۓ�d8�D�3��t��^�����$�_��N���X�5���Ʀ�i�s�����E��E�Yn������e!��}� �6@�l�A�J��Z=�6���ܬ�k#���ߓ4tH/���ʺ?'L?WLP�w3�i'�kD��V�1��.!�;B����Y�M���P���o)�B��^3U��%��\��KP�l�n$�or����S���/>�T�ߕ�.�Qϟ'U6�r��l'Yw�-K�NĩPy��	G��!�>N���O��:1ES�Ĥ"k0�q���MƁ���[r��*�g�M�Z�=�+2�L$7������N���M�`���
Ѕ�4k��1�@��~��L�
�9������U�6����@\&(.��^�ّ=�&��M���x�0��d�G��=��3�25G�;�_7��|��	���Ol����"D�x�e��ٔE��s;
��.�:�=��jpO���ݬw���d������C��1^�� ����2߿�?�l�!;�
�F��y(�A�
�FH��ܨ����>ۙ~66���Gb���l���~-@W�σV�� �v��_� 
�ڳ��
�>#-^��+�w�2g��x!:˗�43� l+��wseFo 3,��4��pA����<6�o.��$B3�yR�q�x壣SIq#��r�c��Oy#�*xg����3��׻Y�	����e�놨�~�n ���St93�/抂ܜ��6¹����G T�;-ya�]������[�v3	K���[����J	H��D���Fά��l+�	��<o�]UWG\����5���"��5�C��4O��c5@�~\-����C���1�p�Fg�����K^fIa65畬b��#�i^�ےݷ����'����n������>�A���U2t�Q�uǰ�����t�M"��r�������ʏ��a���g���2��Z�V����G���}Z>�|1��D���6����s�(����G秎�Z����I)uyHw�]4���9��*��~]/�a�Ԛ���N��$�phhk�Y�š ��,P����ZYoMaa��yM5*5���o�"jK��F��6 �0���$��@	c���B=����uSU�BSO�X����A��~�:cj�]�b�"23SC�|�شvh���<
O����$As)�_�K9
��K-�PL�2-�<k`� Ά�� �ދ�'���mS�D�Ef�d/�i����A��h�©W��(7�C�S��������Ժ�����Y7�B�r� S�`�o\��L�Q��VPf��A�by�y�:��|��8r>j2�M�8�v�镂�6 ]�kd��ە�h�<��I:�^t+�����	ݼ�e:w�����I��zҌP�ߖ˃ˑ�[m�IyB5ȮpK��v�n�5��L�ʾg��|^-��(�?��������K���a�K,:��,�Qd
�e�-5��-KV��G��t��r��1d���<��n��p���:��P!{�ҹ��/����Ua��]d/�{�)��w�F��]��I�1�AG�g[yqw����,��`i}����7�ݨ��T<`����K#�$}�'�c;[�;_Ɯ� l^8��,4G�|��W�5�7��5eHԅ�s2�I|�l�I�����Q�(�[]j`�;\�Iy��<�ߪH�c���ǇF�V�r.��ĖFS�����~����v�A��|����wS܇�����l%���Ft�h��;�SW0C�q�S��g~��"�mϋM������$��e���ec�J��~s����q���r%��ږ��n�L:�~d�X�GxN��j�D�����f�,����k>����Q�y�J`颡���r\��jc,�IC�GLF������8�����G��(��y;e��rr��ȮJJ|�4����8���G3���tX�]A'韸A�?�>B���+������a��aȑ/O0�T�2�ũ���I��I�P��n2E�o��Bq�Z2�L���wP�S�z��4h^�5)�S���yy(<�TL�6�Wyc��Rf~���"5B28ZZ�|����-]���ɻ�恻Zi����3<=x��t�U'ӣݪ�Η�'l�f4!P��c��w��"L�����`Q���e=س��o�a�[I�: �}"��%���/��e�*7h�Ҵ��?�'F�u)��|����i� ���T[:qK��K�`A(�
�<^�H�������X?�Ux�ң~�� 5s��G���Vu�t-�����Z��T���Ŏ�`��k���׺.�d�n=��C����7����?4�,p�c;�a� 	�#�_�@���]Y��"�&,rm�IY��ä$��La���^k$��Y����w�HW��x��s�6�x��F�Ӑ�>Z�R�p[���l��;*��X�`��UcE�8�;k�5�ߚ��!�B����Id��Y��U���(NPz�Ҙ��`��՟�b��\,Y��WK��!b�w^�{f���~9|��l�
�0�핈,�fv��(�`��~BS?��	�����E�Ѡ{X,�,f��=�V����{Ô��x	�?I�q3,�����a�S���s�-�zb2��p_Yb5�^���l!a���2��V`}f�{�� h�0B!��3���z"nu�G��-���8Uh�c�TKY�}3��
�-��R&�f<cN�Y�Gt��G�D�3��>�f�^�}�p9�/�	I�2���7P�ʂ��й*5Ow��0O�8ж;Yʰ�o��+�i��Y��dʋ���V��KFV%�s�R%�2D3�y�|�&�#�Z.:�?�uܢw�t�?�64	�=8���2�:�T�����S���I<�@�e%���n�y���~pTÖ����U��^�똡��%E��;����p<����b�~%�.v\�~$x"����5�;�U�����Qt�
B��;b�&c)���@�ᭁ%wM=�<:�[D�>�.��TI�$#���ڟ��j��E��=����4�7��+&�y�����0}�a��ְ��o��*����lr�M�taN3�S��E����9��O�B8�4#�ek=����l_QA��x��f�!i��z+v�9���}kƃ����iꩃ����[�]¤P��b�;��'Ą���@�!��l�����Wn��2I�~��9�_Z�ĺ�9� �V����l3IS�G���h:���捵gS? {��!#� sI���9�hGi�^����ʟ��9`/�T�8	��� �U(�'��Ն��x��\� ��GW�������M��)C��$@��,H�Q>���cn�Of���#��3�.71?�U�5B�6�%� _�KK#$��k�⵱�m�o��d���Q�!.�m���_�u�ފh�A��^�����Y>tٶ��ke�F�L��3�Z�iF����f��*�h1� }@IpZ(���(�D��y&u�oSH6�������?WK��P)S7$2]}��G��W-��w��/a��K�)�T����Zif/�t߰ݿZS�w���M3z���v婞9-n�X��+�y 8b�C9F!�����ټ*�zh���Y�����W�N��x=\Nh�_h��^���Z����t���"T>Cy����HaG&ua��{|>�t,�F )B�Ǯ��2�������S:2�ϣ�jZ���A�bLY��;hf��'��p���K�����h��!�øB��8W�M:F���&�^�B�
���Y���Ġ+�r�(�0z�`��H��Я���p����Sס�Cl�k�\W]/�X��$D� X���íZ%f��;�{i�Y�����K
�Z�5�vc���PQ]s�`��>�f����M~F�`�}��k+�D�G�+_�]��p����������� z�j�=��Aɓ<-#zZ�Iƫ�h��A�
׬��y{b�3���ݠ)@�E�۪���ը�[n�q�YIU-r�i噔J�ɦ��'���җ��d2B�c��1�L�ȣA���b��2X�N3[�03\��'u$R�1�,��f�q�b^�o���v���=�c�l�;�����$�1��\e�&{��W:�Pb�}�#'��A��TJ»8 �Q�ʐ[�PPV���ыCA��U Azr�`V,����ǯ���d�������=���C�@QE'��p��>A�N2�'ᆺr��z؆@�U�>�^C�����f��N)�����}�aC4^d��ZPƦD�Ўvl"x��@Wm7�^!�>lz"9g�a�c�f�ی���:��'N�s���6J @u���c��v+�M@�	���uh֥q�'����﹊Z��`Ĥ\L�3EYsb��̲
�`����xNgI��޴���{��*�:��	&՜($z��N�������^um�}�k����`���	��CD?݉�2��߆�^��ٷ]Qlv� ��=�C�{/�����3�_�fp��S���LF�w����Y�4Do�J���&}�k$z��^A�V_�� �O���0��2�zF�������|(?��P���[(q�-�)���YVdG�A�$���.��N�� oθ1(;��I��AV���\J{�6�l눳�G�rݻ�_)��W�"��P@�^�^:�B�&j_���`��s��(�߉E�Μ��z��>��O��B(�e�,Ϯ8��`���z��I�P�F�B��������YCV��Qde�����y�YV�%��JI�&q�\�Y.'UI})�-Bb,�IG_�U�új:_��_�#�C C�S�P����P��K����{[°��J�p��$&Cuɵ�|(1��g��y�vgu�Qx��l�"��D����Dd2|x6�^P��+QT�uX����R��륬�`����(�k��X�wN!�͔}�U�zYO6����=�����C9���["܄���^!-����6	�b*�QR������Ԡ��f�J��m��_��C�5�Dj7��B�''���N����/�������&��2K�'{a�C
	l���R��3�����.���}�����Ah�:��B�[.��Wa��Z�m�0���fL�4������l�<����ҁ��_���T��3o���\�5Ϻ�%�	����fۜl:��٫6����.����_M�B�ӝ���"�\Zuu�Z�_�5��a�V-�crw_��g�sެQ���~��~���W�ā;H[NWT�X_�|�F�zDAF� �]9е���sD���L]�7�Yt�9C�W���U���|w��~��z�4Ȱq����0	�#'F�pu�6i搽�c%r�o���:��aMØ�{-u�ʏ.�Ձ�0��6 E���[�
���<��Y�J+t�P���~�<I�5��8(��A2zI�~P��F=��3����Ļ.+�uh&��)/�n,��j�Ց���'���k���A��t�65.c Z�!���4��֤,�jj���1f�b�.�g4H���^�v���̉�è�)��y	��_D�B-F(���H�� $�t[Jɗ.͜��q�/Ã�.c�_di�!�|�{N��j�GI�"J��8I�P+\wx�?��������=ᔴ#k��:�� ���zYr��-���0;.���L�{V2�zYS0�F�U��"�1]��:X[�<�Q�-��lK&t�dMk��Ӷ�{ifAkAĻ���{�w�N��Tɉ�*=}���R w�(�g�v�սw{���fYN�yC<���y�g'��7��!F	�3;7�R�:��riɖ뢤g�̂��(���pʫm��]=�5�t��lr!�19�oں�r�?k���gؿ
uW�J2��&0Y���zc
��F��Mݔ�뜯�J��51��v}�,�vE�E��q��6Z�PG !�M����L��zp�������j��U�F=���d���&�%,���`�E����1��\ Z���J����Wy�o��FV�W�ae?n/4g)0m�Y��K2�����h�M��&���g[������'��<���?��;�w�Wf�=�V?2]6B�`�DG+�N1�.�&���rAI(�ȳQΦ����z�^���佩����:Չ,p�����LƠ��od^΄,㛍YGZ�@��S��qL�a�����D�'Z��Q�/'����MM�(&?�j��U�*N�	��p�OT�o���ʋ95����ZS�'u�h��}��W�Sԥ?g	�|��!!y֠��1�]C6�|'v����df =A�"U�vM�:���X ���	&`�!M�<�RX�f�j��t���L���ϊ�N��$r��u�\X����&�\+�15+1�K�6�N<���ө7u�ٟ�G�F��3k��I�x"-vh�h���"�䑐%nH�Y��Z�5S&���C�{&��f�%��#����]ꫴ�L�h��_�;*!��Ȱ�7O-Y�/�5��{oV*$����Uv��#�B�����(�v����G�����+��ցR����ƒ�p�|�����m"�w�I�_AU��-`�K@X����o�{ݐ��}����{��aJ���W��͋�g(%��BX�3e��t񍬮���
KXZ���j�$�,0���*��2T?�\6h�t��Ĝ��N�M�C��`��E0����A�kG����N�T9}���Y�
0���A�e���|�&5}2o�ã��Q�rtM�Ӭ(����H�;�fC��j3�%��5
0y�5�)�6�nn+W�,&�����H)^u�e��q���\jwM�a������ƉA>���- �l���/�l��?H��T2�܁z#q�ݫ/�ՙRC��&�_�|)8Lh*X��������������8eyu�B���=�
�dhBk3����y#-{%K�j���ͬȯ���U������E�/Id��J=�̖�#�b�ɔ ���{�o���W��1���}��B)ޏK ��I�f-����aΦd'���`}w�t|�~�?��2cs�������l��@5�Cw��*0�NI�����@�}�$Wd��?}:Wä:���> ���gS�8G:TǨ����ޓτEO����Y����Ѹ� �Hi����N8�L��R[�1���R��[����y�`� y��˟]��Y��h���65��V��	�كQph?�6 g�v�Qp�Qzɖ�B|�7�}�`@-v��N�q�$�^�D53t#������ �\�ؒ��I��`��Fk�� 쀙�=�,l0&��e'�)iNn �l56�F�ە���]�Z/b�f;`���Wn���8!��B�K$��^%��=Zr$�Ŷ�Ig���������b��������劶���vu�R
?m��}��k�����T�~��p���Q�x����$�e�na�[�t�6�c/�N.n��'��K�I���#ߖ�C���2�o;<�(PN�i;-Ҏ�N����A�VB�EL��^��_��<����J���$�I��9#�+�y�B��j����%�-�f�ʹ<B�F2���4�n�Z&x�0^p�Q΋�OyOe��e���V�����Prh_"���v��]��yǇ�t����U�.��,M��r��Z]�y���2lO=sZZSL�,|��$ۏ������>�-֣����kG����䒴����mX���<r(�W߼�9�f�ڿ��?*����T��7Ϛ�����_1Qaf |c�ayy�Z�&�x]p4�����k݂P�{��<l1ncr��B�x��o.(5��f�p��Ǎ�3�w-�'���J�����)�P� =k^xs
O8�{�/A4v}b]{M�C���r ����C�607{��Y|����Z�+��9�i��[O�A��(\�U}�Jq�!Zsx�oި�s�hc,���Sĺ?���ѠJ���^��Ĥۢ
ؘ+�/؏E�ِ�Q!�O�0}ށw�=w{�v3c�T�t��L]q+����K��%e�6�Fv#��:�:�R����̱��� ��F�
~{�I��S�ȃe����	޾��Ґ�Ǽp�ȶ��7��`ʳN6��֞��L봹/㠖ˏ�@�IO��?. L!V���Vh�SkB��rs�4���_��^��'�'+�M�1���D5=�@�mO �?�)=��^���ғ�;mj���GKښ��Q�+�����a�p}k��F�i|�ΨڳP������\���}�C�	.��{�1�6�`Z�p�y���p����>�\*U
6Q�Z��ő�f�XG�Aq����To���%�T�f �[�6�����z
�<@�2L�@�ϫ�=]Ȥ�8b��C���+$}�ծ��P45�<���s�6S�wǁ2���`���퉠l5���E��`z���r��a��ey S&X^ҽm�)�}�m���~wa_�v;L�4¼��"	*e~8�!��������*����ZB��]���-�ߔt�W-�|6��`0������#­+тoGW��۲P��@�B�{-R޵�倠��	d2oG�U㉗��}�������QN�܏�H�,.��JE/��-z� ��	cx�t\��γ�-�Xt���@j�2ٴinC'������/����5-/�Q��T\��$x#�b�>B��ě!nT��)���`c���OBu��}��B��*����v��X���ک2O\AJ8vT�8�xNP��׼�s���62�����Ѷ[���F�AzgB7}�c߱W���J�qc�I!NT��l�y�t>ʐ�	m����k���#S�,7��8��M~��7Zx\t�2���ɪ�d��VGF)�t7�X:����/m��g�tAx�lZ�����8�抦���ƥ�9�g96���/��BI�0v�b>��z�/t�c��z�H�N���٧ϵ'���̣� g��8��B]��GC�G�ےb����'������h6s
a��-e�dC�3%�Z��x���[�X��e*�;O�I`���^�e 0�T���ǩW�r������r�O������0�ƀ���΅L�DI�98�^�w���Nꯉ�H�e�>
Hѹ.HW.O��R[���`UAmǴ��x�;L6�E��=����S�__5�/zGA2?�(E<�����A�O�`X��6���A�=��$�5~��>S�������1dT�����4B�e�D�'�SS���{��I+�&���L���S}�]���;�K<�d�Gv�ы�o��/]V�m'I^gF�h�Y�a˖$�}��L��;�A�Ơ�2��}��z#�~���K0y&1�d�(J�����h�t�Q�ǈ��)�B��z��EO�mg�[-AtRVNX,`o�n��	�@���p�`�^�u>�O;~Ƣ~i����S��b��#*#Vp����<����ko}$ŧ�OUl�p�O�!̢C?����QX��[�o�^�yu�Š���R�t�+q���Y�`�Hw���h�s�ͼt��+�F*w�&��{�r{�	t��ea��F+��#Er(��r��+;�ۮ�����1J[
K��:&���������Rţ���ugɋ��W���rj�8J��5q�i��&���Bj�����4��)EP���Q5��lѵ��f�r���C�D�K�N�eӅ�~���w1���煑[^���~��&��9`e�`NE�$��˺�����B�a֗�PRl:�w����P�����[=������z�s�AOp!&�y� ʻ����j����!	%/�q$��Y�18 QT���[�J��<F�D~�� R�"�Hl��D��>�UY�U���b�d c;_.��U;ݟMw�d:��D=w�K���oמ������C�򣚮{�����R&�����'r�� �9��E;[�����<�h��41�,�!r�7eR��@�}�$H#7���о�i�l��g-���q�>ы�=x�)R������u�X&�N�O���<k8Ҹ�TQ�O3�Bhx���m�z�d��#�X汅4V�aW;���G�q�� ��9���>IֽK},X�{%�F��µ����ڋ4��.�j}y�ޜ��1ȉ������)����V�~��9��ۥ8qp�u���jϮ2����3w��#L�8�Ln��n`�'+B���arQ�u𚹾����/����;�.�pI�qpz�dx�|;f��Oݣo���f\C����/�L��^�N���Ŏ�x3�V[Y�$�g	\� �d��@d˧~��z|�m�	�#�Q(�D���3�hKf���Op�=���л�@�nZR��� ��T��6�tsŐ�1$�~Y(���b�U.7ӓ����`-����.��!��D(����C����_ (H���|��Pp!�
��:�G�ż��˺��:�I��V�f���Rp�����]iA��ܾ �wES#���(�en�������g����7g�.T��{�ш��/���8��~��A��5X�U��p�������am���ԇ�Ch�a�o��^���t��S�$P�8��Q>��@ْĨ>�+H~NG�_-K&�H:�>"?�o���H�W�I�>��zx�Lk����!�;G�����s�PQ����ې_Z%��R�� �_��'j�&p�+-�����[y����Vu�N�;kx�fϣ(�����(%��/�=�Y���EY�h�ꑭ �����~�R)��<��+N �4P1�ՙ]�_j���-�+����M��
��Bq;
���enOD�p果�t�$=zd���p^ �IM��<p&��-}�؞,�|��^�t
^~S�C������H%OK��hI0}��R�r��G`*�9��鼀��j�9B{�J�!@X�۬�Wdd�69�j]"�L��ƼiB�Ѓ6�����XT�lP!��be���rBpY\5�1�j;���f��|-3� ���Ġit��~xx3�|�v*-��������~�?��k;BY=H�@.z5I��#V�CxJ�y��Ub���.t;NH7�֥P(�$�F3���ဇ�a�b��m��f=�Q��w�����}���� �i�=�ܼ�v��.rZ�@>��Ge���Q&���u�-�`�ox"�E�,�[C��T܁د���\D��ZR��Ǫ�{EF0���V[�%|��c�[V{Z7� �$��4Ɣ4�b�cjp50��>��3�A�jl->ɔ�՘�_d�/�caYSNK��Wh*�~������#�S���	'rg�bkY^�aLX7k�9׵�r9a��\\��yO����x���8Y3dr�h��6f^8��ĕj���6�GC��L���1hKu�G��P�����
��{�P� ���z��b^.��:u�ˀ���exr�Ή������)#۽ɨ�,�C|R���:��yj~�RD��6��N�R,m�b���)Ƒ��[��ac'��+N�Х^��gR�7�|���i����K���L��?�Mݡ��O�K��6@�=?�
�TƎ$��Dy���ZvL��	�7l|�����A���OC�E����{���Ӝv�6���LXścmQ������DMc.@���F�0/T�NU��F�n'{-Y�u(Y�����ND/��W�%j�Ǽ���r��vV�*�z�ku�)C9)�n���	a�͓�U�:'+'�?ҡy���;��L>���s�W}@��<�J�,���g���y�wU���ټ��U��T��:&�>��fLLF��ok��tH�3���:��%y}|��F{]g؈�|�H�͉UY�����]Ѣ�Z3g'EU�gq� �܂n�/D_����%�M8<�y]U�Ν�^��&W���Ok��x�de�+:�Yk���483x�;��6��`�XO�v��=$1����Q�=�J�X���nq�)!F�ZP���?A�y�գ+�{��9X��-S���K7�ރ�9D㪲�Gp^�������cn��5�
�"��B�Y�(�]�$MT�$�?EGPʹ�$>>4��:��Б3�ʪH��Bn�ޓ����i~�&�\ĜS��� ��:�<\��FB	�ڝߦ@�Y,{��k��4_�\iOڔ^�37e�5ó)#�����UP/_�]�j�֓�B���V��W�>x��p؈~�`�����_X;� �}E���#�kM�|��Y���)�R2�����fF�hG�Ӓ	j�?Q%����c�RFy�:a�p�����r�5�_�=��s|���\3���-bx(^�w����g�`��=�:��f�*=���ӚT��~�
��J������M�T��-xǿ ��*�P�m���G�9�-�R>+@�.��/nOx�c�q�������JQN2z@\P(�%̟����ý�L��3��V��Z�%��%�LE�v�}��-��f��������w�_���ŋU�b|�g����H��K�	؃H�=ݫ�I5U8�K<��Hb���ydU�S�S�����?��ȫT�VN��X�:u��h�tr�8jw�6�����YI�Ot3��0M9�:i�ZEO�ů�;�5z3�3�.
�2&F�!ZerQ~3Hb�)���6�ƅv�ꘅ��2NX!�O:���Jv�[�wf��zM>���ptP��B��0���}=��O ���zLYZ5����Q.�#V;�l���f��G�7SN2δ�`a�Tl3���Uuzo�o��? ����d���ٿ^&	+qx�=+h���#��Ȑ[��$y,]���>��x,�|�&�_Ŋno^��mބ��O)�1�@5�t�Eb����u���;��Lf%c����j�g�R��&����)뮋t�ĚƻmM�� �����2���6,�=U��GH�C;A+ ������rW��6��݈�-�oYa�c����U<�b�Ƨ�O�V=�I��R��ȼ���<tӊ��3R�Gwʃ���$�m���קyz�������[D>z�A�,�0���U�ÀA�z���}�f�}ǭM�)���]��k-��7 n���G��3OR`�NȻ�h3uh`k5��(�ݸ��)���+�B�%+�7��uT7Z��cX��,⿻��Gϼw��t�D�1?	�A�ؒm*.`�i�T��Zѯ6Ĉ;�8{��>���(#��j�׻Y��(+�H�b���r��D�����D��7t��f�R#����8S��$Ś��.��,&D�������yXë����/�,c2�G����:�!r3ޕxD�日(�,�C[<���j=R/*�(	��������q�;�7D��Kh$� y�0	q�f��խd3R�5���>�d&�܉X����fG3|�8�a���_v�m=l�ڞ����h5GҲAa���~����?(�����Q18�����3�S�����v#�J�a����%���F�0����B�,�V�L�cv�C]��f��CB޹��x}ڥi��<f!+^F������6�д���+Cp��0���MW!�^5�����8�U��(ТCd<��YW���8�L�;҇�w�g~J�;:�x����[���R%	�����-��ژ��� r�$��28H)&��,���k5���S�4A�L�&B��Iv���<�(�v2�������".�3�g�i��3�f"��^��!G����&�+�(��C����x�N�z����J	���ˎ�
j$Y� ~te���Þc����N.ص�3��7�)cO�,��5:zR�VV�º�s<����6���ix��O�,�σ�慓44|My��#���M���*�9{�N�6�LR0����k$�-
0z�X�<�:����O��t}���B��-e� �곳�;�{�����
E�D���|T�/2��_s�~�}yM�
�<���i��~�{_x-�����w�R��e�n{� �_��Q�0A�]̺�
����r�
A+�2���@1?�D���x�m���I)zQx�n�T�u�y8
�w�$��L��5|��	
���e�ڷ��4E�S��ʌ��Xh���r��'u��F  �B=4�\��"`���s�<)�ǫ֠ٵ�%[:�cQ�k	a�,-\�x�k"�_��P?0CB:|����e�p:�y^�҅a?І�&�E����at�E��Ə�M����$M(d���Y������JY{7h3�Z�/Ǌӝ
%������M��+�k%�F�[�Xu):ǟ)c�U_D�۞4D�V�5��b���������Aտ�_"�L�;5J;Z�wy=bn�6�y�Y�h�3���V���V��}��`T����3���aS��֤�7��~<��� a�,%�ڬ�װ��N���R���e���0t"(yFu�2jʹm����oE�YP$�H�|�>P�H���h����2Abh�r�r�zo��d3�$ͱ�a�N�Aºi��
���s�=B8܅���M��k�l�d����\~��zIFj;	���7D&+&w�$^�Of<t�W�d�5\x�L�c�%���4�24����#F�6�A�X}q�xS�i��v��s���u<�`����E��\Scr����-0�bg��\&���V���r�����2DA�8�����${�,*3W��N^��iAXl+���]6�1�VΞ���ׄ��ڣ�-"�^��o[@_����Q0�c� ��>�a���z���`��]RS�����[L�������������	A�O>j�� �N����
CQ�LM/��ܙ:��b������	7N���\
y�����B�z@��3!pm�G�n� ��<�1����h9p���f߁F�Aa�8�.�s*����g��[���{��Kt{�2��o�N���J�;#C_���a�Q��E�W��n|썴j�d΅�y��祿 F_�(������l�¾�N³h�����-=+	��+�ǖ?k���X��w<B�d��r�����<�Bx�0Й�6�lα�t��D�� �@�b����n��3�n//6����N��'6؋����Y]c�1�f��N!b�t�y���W��B)(�+u�}�ϩ�x���%�=�_%%�&ք�Th��5�e�FQ3�<�I���v2�	"V8��yS�)�t�B���7�<ݣ�83�����y��gk���N���_>��m!,�7r}���/�=�o�hL+�7~�1��F���G�Νwm�a�P��l;Gk%d�d�\G��\$�u�c����*�}�Cӭ?�9���ϡ����Ol#�hW��<���L������� f��"���]�;,�i��R�F��:XI��*	��=V"�~i�j�m�y��+�N�T�삮S��g{UT���ъ�u�\���Ȳ�Nȯ��{�g����@Ħ��8�\ZH��?b�R8S8Q&��6A����Y���nݧ��_l���������HY�@`��H��I�x�:��Z�aY�t��)?[)Ws�,4q%�A�v.�ƹ~nM�۝�Z%}0Ֆ����xηt���!ӺvS2�)�hJ��+\�P*'���%8�����.��a]���{��&ig4��{���~1�+�M&O��0��*/GRIJ^���f��m�~�&��b
�C�@�H�����!�Xq�5�0>�D<O���cz���R]�{V�N+�!
|'�S������"��Q���%ZWԪ�7?-����
�lUBC�����!�>C��oo�ITi�w�8 t�2���d��`����-|荘J�<(���p�X���8��E����6�x^�M����7�BTX4�D����LϪdx�^y�Q�9|g(��5ʝs<)��p\���������#��E u[��yVL�镎#� X�ei�Q{�p�����xJ��B#	������v�cy��8V�\��u���E��o���. LB(��+�>D�]��g�X��x�uǦ0�B(F��~����@7Х�ċ�(���,\%X&��u�r2n̴A�Üݽs�Y Tx�Xr�v �[���o!Gp*S��0��$W�Z^&��:>6��S�9��b��y�B�v�ǻ�	_+6oqs�K�TM��f9��'� 4p��u�<j�9-Lnf����V.s.Ϛ�j�~��B�|d1qj�4uA�	���2���i;Vz��b�[e
ԅĔO�mul2����p�RP�co�o}����(��(.fnv^O�ti ��
�(EP҄��E��Kv����K"'�Iʈ�o�Պ����'Q&�a��'�r�"��ni��/��!�yN�5�Uz��v��ߑ���Vq2PL�,Z��D&�q�g�=�Ⱦ�d

��Ž-�.n%�����)��+��HZY�4�Ͻ�р&��vw1���1�O�
��р_��=���:�ES�n�E�A�H�|�&ʣ�1B�s