��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:���[�S؞��t�J�{�u��FO���G�+�W��0&��f:]�E�0?�0P� �n��F�P�	m�rU����ߋ�9����j�sa<���{�h�)��0f���.�����!��FY�50��DJ��c>�@�%�������zr����h�i^r}�\�?��5�s�L`*b��"~�y?�m�5��,�H�,q�r6�ZK���~�c�:el�W�xɫ��w����({ ��=��^�莣�X⸽ŪD*5�ĔI���0���=�#,5G�d���I��<l����.�d�O��#�W^Ĭo�^ �]�	+�8ֆ%2k���K��R<��	�佾���\�TR�m�4Ro�[���ZA(����#D9<Z��ւ�!��VQj�a�:]�8,L�r�LW��[X�E��io��y�=$��$]��|<?X<�`�c̦,�#d�&��=�z�$��t�e��qO�X�R�e�H�B�޹8D1�s�2l֐e�a��U)�U�/G�",���A>.�����P�p\�?]ӥ����_ٯ������A|�s���o4�H�]/���q��^���&�Į�'�xw�M�֨A�3�KB��@�F �d�r�1��7P��1WL��w�E�݈��[h�}�1���5�q.Ƴ����(}�/�����������ҹ�x�[~=0uY���Si�b�r{��c��
kÃ�{|� �x�V��b���V�=�����x+�O\�~e��kt���έH���4���:]I�K=�
%&iL�ˊS������@۞j�=(��y�7'�o)}��!�~�BsZ1ifߣ��#��G �^�_Mf � ��������ØRpJ\l��}̒��˫��U:'��M��]wVO5�?k	}�҉����}L���劾A4��1Y�D�����ݾ�Pf�]GI���Jud��N����U�\�N8H�����Į5'4�>g�a��� ��ŻO������Rv��d;��y7?���=���Bz)+�z�x)���ᰢ�k���Eȩݨ�O6�m�VBWco����l�)̛8�n�4R
_�z.�x���4�t�Z��q�);s����`k2�* T�����U��n���ސ�/�WX1�5x�o}g�q�_vS�9�vt�L�v77�� /ݻ?#�y[Ȝ��"��D�F=$�^�U���y�ʡ�&+'Ru��t��!�=��Ho����5I�p�#�o�R�G�D�B�`�Wh{�:����kS�o?�R8�f�b�50�D�O�qqG#:��VӁSҎ���S��ȋ�i��=
Pk�[�}X`���J���Hk������-��ƕ�KF��Fjf��n�|2�LU]R^�"��q].��>N����l{���)��,'�t#�$��ҙ�'!Q��J>�=n)����U�S߈���/+��#��E,o�e Ȍ����G�V������9 ��aO5����h(~��{I"?�G�VL�M�-�T�m��#���`��,�lq�yUT	��̘�֔�P�VK�밪��Ux��J�r=�FeF��MNՄ�,�t��t������/mU�1Vӯ��_�t�qê�����*�D�F�syXX�
��h���qV�U��/ݙ��'��o�]	Ihȏ/��mD���3��*���eءL|�x�G�L��E?y��"���)~DJQ|���'�Ѯ����δ�_ύ=v�2��"�Q�\z�;o�;N P�g*��M�����9�/K(��6�4�/���w�w���F*��9��pz��zb��t`���P�@8=愶�E\ꈧ�C,�[dQ�
��Uv��,�FD�*��V�T�7�EB�� �A���:f}�
)֦������(?�T���i�a0�-t���`����h���OI��L��"���I�'��GQL�ܮ�5z�86oQ�g��B���g���gb�M�@��Z\�dA��?,�� �?./~?��k�������x���C�4�sp$���?x�]Iw;{��X�fN�h��Eg��D���E	�2��ˁr�P{��5:�Fs:j�]6�"��V�
�\�� �i6ꖺB鲛-�.�dm9��Do�-�L�Է���to��(u�|=�|��_0O"�F��^�����0|�K�({�uB����sx�@������ug�p���9`Gx��eU��Ie��䢷��@��-��=4s&��@='U?)�*���A�k�7¢Qp�O�ƞɀ�ʣN����q8�����*����i-#J�8�p>�p�	ȃ�E`9~�m�iVa��X�v趋������K��<t�"ix�w"KV���8N�$?�˾�h	h(��Yэ/t�;�[Mנf�^pcT��vK,�/:٪�;l%^�;��_�VNs��D��V�g�F��6_���sO+Gld��0K\}����1m ?TR��;أĀRc�66���J�VqP���YA6uZ)��ǻL�eW�������n-{�-_�&J}��}����ʡ6�ʞF#g:���0m(H�U����²�Q!��v���Bj2��.o���Ʈ�$�ܗ�3����/�z#��Ȑ�?��lg�N?	��j�]�Ә�m���tW4YwU����iU��x�m,$�ᨱ�_y���N���b�)���Ω��ɟ4�������F�t���Sãk�f���t��1�=M��i�>�6/t&�w�M���o?z?1%��ܠ�4���nA�Q���N~:~F_vm��/�����qW��W�Q�Зxe?�w��������u9�>-�f�*+���m ��|��h����屉���3Ӑ���`B@0�

�]?��;]��aP�(���i;�l��1%��_��k�0�c^�.\�Iu6���݇M�l��W�n�R���FT����(�������	�Oh20��	s��	M+I�Y�Ξ�]���]{�ϐ�]u�a벤`�����[p��k���6�M�t4���]�ME?G@���si?t��M*:"�Awļ�,qbv���u�R�9�k��)x��C��CH��t�4�+V�i�U�e�͜���\5Z��ԋb4!������Q3�Z����JQ���{}��ƈ�⡨���/�X�K
4�\��.��y��LނG��Λ`�Ir�%EO)����o��2�/�Pd���a�z!�!�jg<��C�����=|:�E��5�0q~l�1X���X�h�Sk���G��i�>��-̛�;'?ƻ�u�js�~���P�_c��){7�ǅ*^U�an�h�S��k�׾�������u7��M�.3���l�%�<n	�/�"��
9��pǩ�{�a߷2��s�~�P*�Vͳ��F�.a|ykP	�^��i/3fY�{�ο\����8Q`f��9�i=� L
Q���&t�~Y�ʥ)E�X�� ٙ?z��'��xY�r+ez\u���P�3+p��qhF��kV��X9�yge�"��)e�� �yru�rp�
�>2��K:�x��~װ����H��|liX�Z�`���NehԪ�M�\��R̕
�w�A*Le��G�+�ۈ0[^r�S��}��mla��,��Q]�2��d������.G�M�c����C�@����G�������<]�&m�����"k��Nj���h}~���Zy�s�����Ƭ ĊqNT��x��(]�ƀ�W�lR�&h�wk��o�����ڞm+{o=�me��O����R�U�0�vP ���-�jI�]y�F��86��b�*��q����g�`����[lh=��\7���n��幇�ep�7�?߽�-=|$����
k����7��>�oi�+���<�Q�p��e�:N��HR\) 8\����X����s� ��'�9�$j��զ7���$��J�bWS[�g������WEW�����M��s��a��� �à���g��[�xǩw-�ˍS�q�Q^_��U��w�@��t� �b�
��#ȓ뾥t� J�w5\z��G�F������a��{۹*�� ��5�WIi��mC��=�]������ܹ�~缪x��^]�	:�Ï)�6tr ��X��%���&U�@+��L"�+f��=�!��m��>��;O��ٌ߭'�� E��]����p�#W�ww�e�=S`P�r���;E\�C}���$�6�K������N?��l�-iۓ7d 5=�=t4s�ۉ!>g��t8;�����A�~u@�gɫ�NUP
�{_�M�Ux���w�y��Z�x��^'��u�ȴ��\z�IE�9�`�Ȥ�k�΢��G��X���+�~��6����9o���
��,KD������r7�غ����iS��߰SϾ�j�х���-��0?my�&�&�t�|+9�Q��y���& ��hNY4�%9����S��GF��Ye��$�} z=7"J��@�AN�c��%�9���8f��J��l�MW|O0L}C�{CB�k.(P��I�o�B���0�r�H���Wf_H?�W?Ek�����)E�#�P�ؒO��[��Z�����t�B�:�h�T�����W�;uP��ɂ�)����𽛞K@M���Z��\�s���<�ԁ"2KB�	�y=[���E����Lp&lC?ү��k��ƲkHB�N<��U�0$5A��*uw���o�b:W���9N��B�!�rD\t�7�ӏ1����8V[�6�u��#��ieg�� ���Aw�S /��M%�JG��N��L�E7�௴j3��j�?�V�'t)�/ǚAqɡ���W�����v��;�1�������1���&�-sx5ַi���7���G=�FGv���m�"�ef�p�� �#A���OdZVY^U�^�k��O��:�s�A*��f�5=[�BB��=�ڟ��mƫ�wO���;C ��\7���g�gz��,�U��v�;w�b8NE|}ğ����� ?�٥C��k�C
1�~k��
��N.�t���x�̬
�Px��A_�Ȃ2�إ�	��E��g�v�U�t9p\1m)����\����cI�W^��v��C�%jf
%[� �))�v��9��2ܼe���O�sj+�P�c�N�z��!$�,hW�s�*����7��ᨃ�C�m���{?�\by��� ơ���ٞZjx���7�I^�7R|n�b�� ?Q[9�[�X��c�ƈ/���,���M��x��
����D�Z�ZoS%����XXH�.5���tW'I	�'2�UMܷ�U@��+]s`GІ�K��i*����'�δ�������1V�eLf��#�M,l��yщ��n��_L>c�g"4T��K�(	�u:@
�X]���M�� ��-rp�Z����9�R��y�d�􁬖�]]b�A�)���jV����x��<�˶0�����;5ќ�Mf"�A�}(��L����Fm�d �E���a�5��­�&X��i����<���U:��0���ʘ�6T��{N��Z��kp#i�ƃ!��c�a|a�*����3� �}�o���$�~��;^�,���Ns��]4���u��ޞ���2h�v�c"P�O�;{9L�B-c�����Ӡ�=�<��=�*�s9�N؃
����Ąz3rm5,�o�|Q?*��_����(8b�&LdnҔe*]�ͦ��.�m�I�{.�@0�e����O�����H"7��킒��^;�ϕ;�?'��Љ����I2�=�LG�	�Ŧ�K�r�88>$^����~&�t'���osѝ�XqGע���`�)km~����`���{L�DN��]�oέ0��ny�e�r7���`mي�"��L������vF��{y)�~_�Rm�O�)�D�Z�Rz�Ч�<d��U�v�n�&I��9��Yr������Y�J%z�5WT���dv�-� t��e�E\fŨ���!�Ar�c���227�O�����C�4�v�Ò��҂<`L,ƟHw�?P��!u�ym��A�>���%C��>I6^�G�t�_����S ����s�F\�]��,Q��J�����\|?��{h�O{�D�G�z�k�>�;9�k�2>l���(d�x�,r�CЮ`n�MUfM�wz$ ]A�{f�}ʳ�z��i������Ɯ3���Zl�K��v�����x��{Q�Z��*?������p�h���@��\��Fbb���$�j��w=�]�	��F���֍���a]f[N���� ]i�봠t�������)����+��Y�M֣�zdq�u�v�1�i3�C�����K�g"�m@���}F��jj}Of6ٳ�U$V[��)��۝��2˖E�.��3[��Q]��G� ) 6��p[(ȩ��
7��̧�tQ/;5z�H)hh���Μ$�e-ddQ���26*SD*�Y�=Fl4j�:�o��z��}���YU�������G�6�6����R� ��b5�4�ƦR)E{���	ᦢ�6��Ow"iG��Ӷ�aAx,#l*N�c`\�@��'��	}��h6g@@�/Fal����[?z�����c����_�+".�ށ�]^B� �)PIr�uQp��}�l�<�/�.��@|�#�Vw	<Ǯ	=>Kk�v$�֝X���𒳈�Η�R5d�B �H�Iltw�_���a=�oFl��a|&�̑������S��)O�0��v�8Y��eZ���7e��~v���gkG$�#D��#bo�B�B�����x��k@����Mt�xE�$Oٛ�[�����(>JUҚ統*��1�DOc��s̮#3o�Cj���A����� �v�K�#���/����wC*v�З��nꔖ�E��FNC=P��th��y��QĔsv�������0'!�=��^P�6jZ�3?�cPWȅ�$:`q�[�n�(���3F3��ŢK�A��R��)%T�t�%6!E/N"�s�Idz)���� fd����44tL����)������!O��>�1f�l��]�IK�s���O��� ��(1��@ʞO$��P�4]���k]�G�DQ
1��}�9�H��93xƁp��.=���J�~���&}3l�	A�D:��믚�#]\-�id�1
������\��C�.Ѣݷ�] ~V#��pX7�B�6��R�DZ?��a��D4J������#�����?�5���R���j�#�[A��z��.K���Y�v�?m+���<�DO� ��H0b���|Hb��{���y��6���`��k`hc�ڑ3�!DuMg}�����%I����Zy��� ';� 5��)ح���&ֿg}{f�̫,T�ڍaӔj���G�݋_��Ӆ;����	;��$$���g��l�!NON������V�ǝ\M₥]� /��-�A�r��NY����H�� qϔ�v�,fe'w�/u��-!N�!mh8ځ>�L�}�%PcD<�);�]��ݡ���1�SH5��S��N�������8��`�wn�k���bwō�����u>[��tw݈�<�!a3b��ɕS�J�6�II�WK_g�hYR�L�� �kQk/p�"9���i�_=Q� =��*�Xk���9�s��:(�v�㾻-;�3k[�YF{
sPՀS"�?�X����7 ��8 AR�)�K��)i97}�!����HG�5Jɮ2��c	���L��-�c�Ј��a�1��:�%��d�&����u����/*�M_��2~ٹf2��4�����V�M��T�f�E-5���K�L3�:�������8B[|�5��K���Bٜ�٨�}��s�;��ٳ�|O���?ةB�	a����i�\�NJ�%��0�j\'�Ade��/�@>=��k�f���y�g�̘�':ގe����\�B��̪ ��=��m�Qa������V�|�<$q#U��)�V@`a)�h�w��Te{�Y��D�Hj��f���^���X����Ř&��o,�ې��:(��(�؋�$������5϶уA^Q;*��S0�^�"F�[q��kR�����3>����`LYh��â��e�\w-�C
e�+���B��r��vtz��S�0b&n���#q����#�^����If���A��ś�#���fl���Qn�O\�yU���IMɘ�y`\ٯ_o�j�q��̒��76���?]��њ��v��r����{:��e�St)d�@�;�݊���縘E�*OZ��'��4����5��%�c*Bz!���2����T$�j煟!*��,M'��X�HĒ��q���ѵ⁥��
BBƈ#������6�Cnk�U��G��J��o)��T�p��H0����|~�Uco7�6n�$3Z�C/Jԗ,@/ /bV�cFؓAZV�2�!�֩�d�������[.�]��Ż���K��.UQ��h�T搤�,�J���}���������#,,��L�p,޸��;(0r*#�b�Qu]Eqmcp?�G6�j���F�۶EXE�'p����;И�hy���7[5����E�����v�>P��#�����%Wq���&��Ϗ�N�����>��@Z,V��3	}�����z+�#���߰5��r�Ϲ�<�6C�L�n�3S-���Yst��h
a2���e����fJ&?�˵�2���˪ |�J�\�>�� �h$H�%e�R>e��S�`����5���9H.?DB.ʛuv|�{��kQ�*��C�{4زbqh�
����6i�og@�Oހ����{��9^��1���wgo'-�:s�f����#qlde���]QƓ���ιK��`�Z ���8�{⪍p�_��!�C&���-���CLRwuZ��??�����G��.B2�F����`b��[��P@�(���˄X�/.�d�q���1���U,�ϗ��Ӊ���~ #�(��!D�c�he2�G5u!C�c���Pj�($�N-�p+ہ�3S�L�]�=
oCHɀ����jw��026�_��g�iR},(])��h�P����)w1��͊�X� �+L��1�A׭���Po�Q���*}P,����jBvw>7�I,��Z�t��vg�{L�ca����b-8`���!������y���vs�/=(��гS�;��B�~[���Q����猵:�H�b�.�[�Z2b
󂇶1����f�|�~�]w<��k�oS>RJ�9�@c�\-B%4��¾��<S]��/<�%��ڥ"Q)����ynL�hg������T���3r���9�oFNH�s���FR�ͼQ�&g��蜊n��u��ft�b5U��t�
���`��V�$��a��].=	�S�P�6��o�s�0O׮�]�낓�k%�rl�=��4,�����Ԇ��l��C��E%<"��`D+��"�����&�
͆O&�K��A���H�?���;�S�l�l��gV�Ij�YH{�@n������Q��*6� ����CzhʁBI��Vck�LD���R/����ݭ�Rέ����ҟ��,.����>}���1���c�Ґ�0?V�p�r>�b��oݔ,����R���'^*jy�Xg����׋��-8r7 9��]��wQbC��K����+?T����͝����%�f���/�r�^#vb\�'Ij�z���L�	h:h�Z���Q678x�f1�F���&NM��Z�KkΣR,[�YL>ߌ.������5uH�8N&o�����G�o��@nf�*eU��v|R����;�02��\i�nQ�!�@}i���;c,��ըI0��$^fk�-��夘��'�\�¬,ʵzI����a@��Г��@�ƻ{�>Er�^zS/K܋�ɜ���y���mBw�lJ���j�'`�\`�Y��=�A�|j��#��)<ylLH��9x#�|��q>Ӗ$���6���7�k[GS$��	��m��9YYE����<���Y6Y����
MV�Ř߻۟��Yr|��5��e7�Dl>w��J���tX���O�}�=EmA��|�s�a�wnt���3?ϖ� \H��M͸2S16�����n����S�0��m����Y��UCE9�"#�V�f�&����(o�z��na�]7��`j�_�c�-�9i���9��j���N�y{�/X�K7���?�_����N��;U���������ߜf�G}Ϸ�!&X�0�"�+?�S��s�*~��� �Ml������w s �n��-�����2M����+��x:
R8�r	��QX&�Ā�?@���
�G�,2)�a/�j�5�0�+j�����t�XL6!j\���1�[�4D�w
	�г��p,x���D��1�?޿�b�6��,y��w�cޝeJ���6N=o����B�QC-�jj�x,��x��S�R���`���Qr����x�Iƭ�_M���2�[q�LB�����ة#5�T��U�V��#<:���x��,��6���Y��B�_z���ho����T���*�� ً7����=�O�i��n�|�e���e�I���/�СS˚���v�D��Zf�,�̉)99.���<􁿺t_�u!�G&��8Im�	���