��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V�K�=Yn����H�oe+E\T��F]��f�<���OOl֙�7��-�Yw({��e\��Q!��|@Z�p�F��R�]�}ghN�>S���Ʉ;m)�OI�� ��N
1N����S9�r
�ab���JA]����������̻y.)��B�o]锴�."�IY���ǳ"�IƦ�
�-ۥ��3W�J_1��|�>��"��j��0��Mt��3����}ʖhb����E{Ӵ��wO����R p%�5!VD�2<IZ�tK[�� �^S�tI�w��Ȩ�p�W�џ�&�m�spY�׮JjfD�����w�v���s�,�Ƽ\{^?JQeЌ(Wv=����wY�1�w����G4@i֩j}'�(2�\i�Y��έ�tjw�����B���g�L0o
h��]TN��q�l��O�7��h�JK����"�ԜX-��|�	Z��G���u�� ��2�yC]�Gy�ع��P����k�����v��=��2�́jR� [<��ɭ���&|�d�l1������k���_�;x�oy��UD�n%Ӧ c�a��0[�oE��WQ��E��N6T~(��<(�%%Px�M(���*��\�����8D��=��[�0˺��)���6�����Db��9 �X�ᜰ�T]�K�n=��<O�M�f��ї��;����r^������ �U0_0s&=S�����׶�����K��U��a��7԰^J�Q�hw�<��є[,EP�l�@W��z{�e�q���Kpb�:V#��S�N8˴�ٟPQK�9�i�uو:�b��e����Ul擵5AB��A���A�'[�*�X8��ˡ��d�e���f���3��
�e9��J&������
~8
��K���P��yAo��&�G%r��J��[ǳ�c��#gJ3j����X�)�81���?��_��c�k�������[��X�_(�|��C��%�d1�[�����H{���:��F#�O����z�ȯ��˄H��g���u<?�şC��jDB�W3](6�S2gf���ӌK�ɟ��W#�iR�|{�qݗzbM0馼Y��-	W��������h��B Nёg�,�CjT���\���b�Bl���LVޮ=���)o�H͕[~��*<�!���5PX�0�k*x�^(�D|J0��L<��ei�3�H���8nڡ�^���R�