��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:���[�S�3��s�?�P���n
�Ә��\Q�^�ĘץR�Dx+�Գew4t1��i�#���{Mz��u��'�Yc���f�( W���+�����8޺���^lg��WԞV���ߙ��⁤�z8�M�M���>8�r�{Oӆ.���Jv�����7	!Uu�IF�1
Fy�P9�)�	����`7�/ү��ZR���;��;YcgJ�����s+U��K�ќ_ji-�P�[��G�k8�1j��zpS�fG�b�~%�F?D*���k>�2� ��}m4.H��s:�f�fO�9�f��������E��$�f �kmq��a���U�պB�U3��ev�*���,���w<֧P�He�9�@a�l7D���]��F>�왙�����u�����Tgw ��%�ۖL���
�n��Y��]�`ң��/�b��UA?�mW�ɦ�sP��O�a����G�"�:sr�ë�)uĐr���U�]�XL���c��"g�Y^�gg� Qy��\F���4�9m�d���4Nڑ���s/�(P���AÑM�:;�x
LD�~~d���\�Y�� ��˽��ez���$�|E������� h��e&���j-64~S�'�\]�� r'b�((x{�H]Gy������X|�\����8��,)f�܋������iL�?D�n 'zTi�,�ы;G�n�?+Me�_���u�� �**0�5��i�+�8��FO��68Ѽ`Su�st���@'߱{k��e�R�%���o"������A�f�9Z~2�U�����q0���N��Z�9Q�9�ۧqT��mx�Ҧ�M�d�v�B{�'O;ٞ`SL�|Ƴ�c-���a�y#95&>�&�ys$E���@�T�v��׻IIO�	�������?�=��5z��60�&���r�2ͨ~�o@|O�7����zgHs��Fr�szT?�}�I�!��e��G�ǕT;�4�r���g�r*R>�pq�P��L)L�ewh��H����鿘}I��Qʋ+��n#���$��O�b���?��Y��3�1ˋX	�61��q�Mdn���#fa^HL��M@{��-�>T%�'�5���X˺��pn�r�R5���&xK���]߁�-�YsG`	b+3K�V��MUi��2"k
�`�:#�p: T��K�m>�����+L�G- ��{�|�bo��u�Όo����t����}g�K����L����tN�̈���Ş�׈_r�צ�At�,Tʞ7?�K���[���pN"�&`����=F��V�������"�N��#����R
?| �9�x@?+�$�@�:��튟F4"P��M�סU܆��P�!hI%�QV�.���d\��6�h�4�:ý�N8�
@�K����p}+�p��S1�`��\� <-�I9[{�Q��ţ��u�8��l��h ��� ۈA��s愡�h�E:M�=q1��l�����tR�y����7�Z~Ӭ��I`'���c>���0��0&֋��5ѣݠ
�߷��:���U�D�gmg�o����r���F4���-6�j#0�b^��L��K�1�������8���-�b	����S��=��I�{,�2⋟n=G��Qx�gwtWVw��j�R��WQ�Ȝ�J�䌔�J�Y	����9��46.��x��X7`0K0��8���5!�|t��S>�2�2yW�9���dP�ffMˉ�+`�
����f�b�m/zs���mE@d��=�i,��6�4���¾�bi{�����f�{�%���Y�)s#}�0>�(��Y=��!��y΋g2�P���9F�����q髹�� ��U���R� B Uw�m����y}N6Uّ4c=�:cc��.�K>�*�z�h�͚ȟI�{�$�I�U'��!��V�~�&�����|�O�_�7G��ĿUe"��R�S��H#���BG	l�z()�a��#�ޕ(�D����[�T�n�@n����戳ILHKߐcf*�an��pY�RdW���Ta,�0N��ݠ��*�E����ŉ���{*����{���]o&��r������O#����Ye�'ޱ5~��7���\SN��姜�
9����i��?�"��rx?SNMߙeCN�����F���5��kPn�/ёlS5ml!>J �ۃ��B=@��=�n�8�NE�og��*��t5Ӝ���~vpw�n�����iݟ�����H1v=���T��Yy%���$ź���m��|��v��P�~^���k	C������>Lފ��l�ۅ�G�(#@e:t�j����״[��
���C:`1�N�"x]�e��ķ>��.x8�i��,xn�к�$M��E2l�J�.�#Ihh�B�_R��.��tU@��'=cF]s����p��b��:��nѵ���o�W���gN�n�=�#��j�� Č�}�ᔻi���$����듉g@$D�n���Y�
qS�#�� �&�İa@A��� ������t�Q���6�%����7�h���<�?�_������f�Q;���\Ɋ��Ώ������x�#�1.�\��Z��xP.��}��</{J���Ω<��X����m�i���q~2�e�֢��V�R�����$=������k[��<m+�W��� ���	}Z�8.��*�UxT�n!෺� ���Po+�~BU3D�1�(��*��$�;o��>[�?��.K��y���k}=(���j��5��k����lw=�<*_ ���R�.^'���2��B��3�}>9^)�k�/��G�8O/j�|��T'<��f[u��G��&��y��G�Ԁ�i};wl/��O�l���s�
*ݱB�$C�c��o�zK�8��:���y<X���l?d��� ����g�vx�P�|AD�>�ͻs߫�ѧ6����J���O��NOc�*7nt�V?Lp~�ǜ�a=1|�e�o��8혉a���@��O��"� �q(�l`z�,F�O�W�����d2�G���n�J���D�M���>,��q��u'����7}%=�Z�~na��1���m7��8��M�[`c����sBq��*�*	�M�hw�jD���B#���^U�Z}w�m)�R3Ҽ��rv�i5��71����A�!�!k���	�`�/�D�s0P!�ˋ�n��Y�퉨���N,Ǧ��+��-��ץ13�<�*o��"{��]���-"�{O��b2e����܃A�!0grnF�}�����v{K֖�/��HZ_
�w���U�ܱ�@�Wd�cZ ���j6�����IŽU�`Z}ꢆ`	�^��g99������F�����Vc+<k�K�ܬ<��h�H���V�,_�	��b�X�4�(E��ff�h�"uA�`�^w�w+��sC��C	��K�>��كO�I��麖9�T��6D\���g}lP��xκJ����K�3M��؃<�e�;mI�;B�Z6Ĵ��������O0��p��|ց��'vB\��fL�$�ޗ>#�p'kp� �g8+��#?V<�B�PA"�'�߂Jh��E���fo��+ ����>m~E�.�I��`=�	!@6^��6�2.�����~+�we,gr�#�0K\�����%苹r�N+���h/��߀���Y|0��~rj�tF3��;�K��v��#��m�wʿ`ّ�c_O�u��':����К-�R�����sp�2Ct�;���P6]}�4���ì�7�C����D�q\}�i�����a����2����}*~/'���"*�>��TP���k�K�,�x���RF�`7_4����RG�"28� K�tO�����=�����@{@���{��������p��Q�T)�3��{5o���:�`�-����Aֳ�|���X ݆�
���,A�^ʞ�ѻ	K/)Pr�
b�B�$a1I;M��Z]5J� ��#�eL=v`d�XB��;��y�(�``U+�]�E���XG���T!��N�Z�+�8��0�ڛ�6�[.m󊒟[e� 5Z�'�ec-�1�qS�DN��Ey#(芋O�M����1H������H���|[��D�<������DG���u\���7d5͡Q\+���R�&TŢl>tP�V�I�p���b���$�Phx/�'�WV��V��� �<�H��'L�TqJ�X�y"��g~o��slkH��`���[7�
����d���&�R���\"֔D�7_,W��غg��Y4��Н��):�g�������H�,�ik��]V�3P�͜������.Aс�2��f�h��Oi��uϥ����o2!9\�y��zaU)�?;���(F��,�#Ď��S�A)��BlI��#��L�z�lm٩����[��YoLP^@�����pr7�F���!/嵪��Sy�V6�Ovy��\ɿ#��~,�JC�뒘�y#Zǁb8}���\� �B���q�b�t�+%��὿{N.�Ѥ��X�H���J:@nr={�;���;��:ϫVѪ���l���5�Gw�h��E����w�@�ɣ�W=�O�����'�Y(�m1����5��\�t��4��Ċi�Q�M�a�_j�R��f� T齠ȰD�
�|n6Dx��(�h���ԟ��
;�1۴��X�^�)��oV�;�& l)��_$�!�,!�2P>��N�|⾭�۩~b�拮��H�-b��o�`��x`6z;u����W!yfb�:`�2^n�$rF�	)�њ���0uZ�C�] ���V��vJ8J>��XG��WD�����\�	��*����d�y��v{���C��Y>����w����ٌ�<_�p���l��W�dX�E* X��ct~@	����W_�ɕ���tk4$�
�h֐j��t9Lg���\%+7��h����|��!�4�`l���Ѧ�'��/��Cc�����)ˬ9�*dU/�,M�.���!������jf�a}$d~&���IL�8�r�[BO������ǝ׌�Lob�g�[��*ߧ�0ɝ���!~�+B'Y0e�^qY��W���kR�P�+\���7UD#����)�Đ�|&�F�٭�T�{�g0�'����q4񂉛ϧB����yӰ��˻e�?Ѭ�^��w�SS蟸�"%��^��@c��̠mU=X�ʺ�f���}Qi^��?��c�!�$��ti�OW��9��@�\ �!�Й�u�=��\'Z$K�#�%��n��Q��P�y�j5� `/��ؗ"��E�1t束������4�4�����]z#�d����2�9}Y��Z�7�#�U�b�KˍS$�5[
��'dY�p:Qv�jw[���<g���T��R��ƌ�;%j�w}Zf�=�zQE��Z@��i�"���/0c�Y8�s2���m5�ʐe3����okεO�r��-������f���ؽ�ݖ�9�J��/c�8����?��2�����3�a���s5&ʸ���nB`����:C�M���M�:d��$�-�i�X��K�D�T�.r����g:v�����8
UY|�r�DDj�Z�;�E������*+gX�4� �8�Χ-�zڡ�Rc8���	g4Uu���n�7�O���p������M2J�W�z�����>>��9�?TX���Xj�_t�[4�r��C�^��~��i=!܂3���&���T�����F���[_�R)@zDl�� ���nC��$ɨ�r0S���(Uğ�����W,�v!�U�@��xj���jeMHנV���>T���9�����,~�T ����)X����9/�y���i���n�ɵPýs��$v1��tT���az5eYgjx}�ˤOb�-�燂��]̲oFݘk����OC�D��W01��<���-E�����E[`2������c��&�(Yo�֕�`X~���7�z��_�O�V���{^�Xi�W�-�&�+����(����Z�|k�ܲ��M�u�,�A��z	K�A�s��/�=f� �&/��]ߩ����`����S�Xa���N~Ф�8k�E��6��b7�+[K
pokțF���_>v5,� a0��1��y����}D�-!���nY_���[C�Q�cLB=�$����$Nϔ�q����d���j�7vm��7:�sՌR���%N�n�u�Nvrg�ऋUB��D�
7U~d�EP�������j�����5"���}@�U>!S?@�����*ú�@�� ��6'�4�m�,ߗ"���PF	D�UR���BK[�kkR��uLi������������6��=�^D�N1X�*��E�f�O2���JP��yX�ب�ԘԷ��Az���*�R3 q��<�.1
+�I�Բ`��U)ʍ�_gN4�]��K�k�.����4G�� J�^IʘDT�'g'>D�!��%��
���������v�~Qؓ8+���Yؕ�`�ٌ�]��	�-K��F1��X�2{���31M��P����������j$���
�ZqJ�S�L IR��cU8Փh���W3&m;#�������F4n�g��A����2h�{b�N�����ٚAFCU1Nlq�����i�Zz�kJt������g�D�=񁓹<�"��:h-������§��E,n$�%�`'��1�0@���2�ׂs�X�˧�K\�0�g)�Ȅ��[0Aˊy��x�y�i����cÜ��
�F�;�J� �tKi�ȡ�֝�y�4���ٺ,�1V���_��Y�&12;�K�Ƈ�I�����1� n��i�ң$c��,�,Im��� �w ����s�
��s?]*8O����M���.�ۤ�ه'R�Jc÷�c�y�襣5f�6����S���X!6�vq��� �C�r),�ۛ!\��j*��C�S
���8ΰs4-C�\F
]V��l�˸'��?�]��Yw��KB5�N'N�]TĭP�s��� �b�P��T!g����/��4Xb�t�9���$�u��á�m?v2�v@������%j�i4�t�̈́栱�W��x���l�)9ξ1
.u<��M�j��(�<�5�x�aT�L���/k�_��2�M���.Z�����`���d$4]�9>m���|��$�6҇p"5��~�i wN3{6���x[ze�ܗ���R�9>�k�~���Mq��=Qz{�0�"J����׈���|��1�$��1��x�lI�o�K\Y��J���n��@�L�!��a�<����M�ir�	�������!:�4s����A�&(�/~�&�P2x�f	��*��A�D��M�T�ˇV�[���fɦ{r����߀~ۍ�*�lO@;ᔡz��t�6�kpĈ>����DG�aD�S�NiZ���$RD�a74<�|Y&�P�wP��2|� �*�}���u٫��s�T/}���_w����=�	P��6R0���Nг�@��}z��4��Xg}P��k8��K'�c��(���2�VۼMQ%��# ���7L��_��l&|�Nn';�  ���� ��!�ړ�,�����@��M���R�����.�G�{�g:���7�!����ʎ��qs��;����
��W˚酕��]�&�n♒��R��/�=�꒰ �d. AbO��B�r~��a�=6ĸR����ٜf���D�ɓ���+V�8��a\!ۙk�����P���	�'����W��3����uY3{3��<���j�:�^��Z�i=���C���:�f�{.��3���^���E ��R�^%AA�RR�2P�f��%����A�T�7�Դ��M���6#i���7�4�xm�6�H�s�_q�HRCZ���)=�d�5$�t�1��Tp>���K��*>s��B���=�yA�l�<���p�T���#@ROy�
�|��v�ɟ�/����6���́|�4���2���^�^9n%�-�k�#��
hCK����P	��dE���ߌi�����_�����"��e�M�Y|��Sw$��C
�@�R��$6n
��O�N��5�^���DU�(����Mq�	�[q.�5���U����t�묛���=}Q��j(<�𿖜pRO����U� l�N��G<��W�R���s%� \Z�W#`�n�.5�J|���T��<�(��D靶.L�`AĬ
�#�=N���t�������v#YH>ćG�	�7�e.=�W
v��!��"mt��W��Ӽ���e .��}��Ի)����%w����[+Y��M �;�P�lB0��Os�Jȣ�-גǖUݿ-��ۑJ�@�bB2���{�6@K,��$=_��5�|������#+����#�7��R1�-FQ�2ڽl#S��h�r��9U��Yɛ��:(S��1����9j�N4��uOSᚒm9¥�6���E�|4���3�F����É
ބ18&M"/U8m��)|?k���-톸�����X������عl���r4ޠ�!�J,R9��M�X��q�_�ߠ�yRe���nL�[a�����h;�-b�5�eU.�4�q�x:�(k����`� ����I�0ڗ7H�� O%c���'�J���a2��/�phc��q&�ơ�Mbؿ;Ţ5�u#�.F�/�5�okN�� ���8�>d��N�Bdw�};�Y����m?u�|ܺ���.�z��9�*�`��M�1RV~M1�i�o���p�	�N:�i2h��G�}϶�$9?���%%�,z����׺W�R4���t�XGԪ�
�\��z�0������׃��t�7���FO}���?�]������j�-7n�w�Q5-ly���������D����W��vH9�*��|2a�����e�*^g��s�>�$�b]xI�}0}4��6�s\1�.�$LE�Ut8�T��誘�� 8���'�Vc����-�G������t@����.;�}9ҟJ��0h���4�=IK4���Mշl�>Q�|up���*+uNXL���s��.��S��Ou%:��CB�H�o̯~J�ڷ�h��Ⱥ��!F���q.�*�8���� �Ս�CDo�3NOÎV��搹'J_]�K�9�_d�K3q�dK���Q��(8�P}��n�*����յ	���PP�����Y0��HD� ؙ��"�(��1��Iܓ���=�6�<��,w-�%�E٤�"~����qU3zJe�´G�?/u�-��ݨ�5���������k0��6�&�R�7lCsjX<�_9.4 ╡��n�C!7'�a��ړL[+��4s�~*p�TX��;�P�u���"����^�P�|M����	!Ta�G�Yav遝�=1ų�hׅx�  �l��_`������ֿ8�.Q�&Y�S��l�M��p�	J���Nl�;�,��bҁ2k�cif0Әu� y�{���E�n�zg�M�x_-�u<���r��\�scYS��쿵u�I$i"�kD�l��ƭ>���'�b��am��j�&}�	anh!�p�n��E�(̴@�ճ� ��0��[����O��^���o^qyE��| T2*mp�)�6�YU~0����!���솪����i�r�L���^Åq���A���󁨘v���pl���G�[;�$��%�vX�p��l�Kd+�<��a1~��ɷ�)B�٢��F�vϙ�
X��*8�w��H��[���\z�E�o�n��k����� 2��&���X\���J�1�K�J̉X�I+��T���W�/s�Ɋ�΀?�=��Щ��Cb3�mN�:�8^�p��u5�&H
_��;B^iՄtg@tU#�5��5-��ސ�o@^�e�{��O��