��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�U�v"�5���rLRU����{���8,�g�1*��)�����Vh�4���[*$�v��_Hn7��,=��R3O9��#��2@v��H�(Q����nQN�%�B�G�>60�ӥe�:g^.?����6.�IKS�ױ{⮿��p�pË��_�&���!4b��[0��E&|�:�N�2�8�^��8�ё'/ދ�y1�ʌ�%�/�&#@��6��W��P6�o+�-�+��L�R�Mz>G)�)�U	� �7�1������BV��ı�b�)e@���ES7��������k�F}������r�`z��:>�x��]���� G��{Φu//xb5�>�j����^@��'r��WFy�{˾����{Wtњ�&k�fn٬��ߗ�'Yhjp2Sm(r�iVf+�O@.f�pe�F�K�=Ŏ4�tbK7��ܺ�3��1ɧ�*��T�Rc=�d�{Ș�%�����dR�	���I�:����͊���x�K��ZE�<��$O��#r9f[�5���t����,{�c3S:.�ø��7�i,K$(B������z�0�Њ�5�7�)D����FJw����Z��<����g����~�y�ғ�}��U8�Q{��S%������V3!A�����,�l�
UF86�)R�@���\Y6�gO������d��*l��
�8�o;yku.����l+��[6�t{�K���Q�Qg9�i6}Uˈ�=�/@wt�$��~K-���eL���,^媢"�O������~.l�^	¯�e�t��C���%y\�E������u�����章�����dJ^��'0�=�n�o�\�7�d|Ѐ�}S��"������{1��1O��*N��gT���ͅ憘����v�TE�5���@�8�B�$fr�}8r��zR"RhD$�0ߘ��1�m���%�P�l�t/�^�H��s��_B.��n@Wh�8�7�,1�mԽ8�k�V����I���Y��qզ!��6�������{zs)r���VH"�� C4��x�8
��4Cww"�)�����nx[�}�I<����1���M�B��'��א�d!g�� w��'zY�H��bCn�`��#�Q�>:i����R�gM��k<�F�r���U�>5��Ji��߳��r�LI���$;l��Xzj!����_����A%;��\�w��ﻯ=R�H"�M�Z���)���?�3�Z#�7��1 ߼�ԗ��D�4����}^1�P�c�a��l��מr19Jw�Z�s~%���C�n;�ʝ��╒|��
�q���C����m���b�V��,'��Ww�;8�_W�YT{.yR:{'�å'��i����}���te�T��IK�%���K��7��ϗ7�T� ���A<��[�d"�+C3���Y��g"!4q5lh�ԯh	#�7���x��G2!�'lP}�w���W�
�����~ j�h#��-�%��]���o�%�9u<J�Ov�T�_��A �yF���U��]�m!��ub��� ���4
����念��G<���MO:ODY
OY�#�1�fR�.�i?_���1�\W|�Zh���x��ߩ�yu ������j"jO��?$kд��;�M�99̌�@��̌1QPLN�WA�N��3���i�h]��Z�C7Os�����ri�%�ȷ��h*?�B���L~e=)�����:�n��<yL@�fX��i�+�UD����շ9W߁j.l��T�[����:����'�fBB 03���D�з$�0A!�>�;?=�b���\E���1үV������<D����	j��A�����q�Sao���������r�w����B�9�3�Ha�Y�^��ZԉfPY�ž>Ů/e�1I�yx[�[Yo���r�\�����?Ԟ����'�G\"�-�P��*1\����N{n��E'�[u�A��{����c(��lY̬ª�#��8	�B|�5�Fe��&+�2�;��#Mv8[ʰ��y����r������/�l� }M��VW�2^.F���t�X?"o�3o�z�1F�!7���h6?�q�ԛ���5��K>ct9T�mA���,�Y�,��^�14��p�� o�a2 �TG��Y�8�SX�.ѳW����� ��&����.���\��iB+U�0A���L�4>{/
�����F���}N1�(MY�J����`�E�ǁPU��>�q�� �V+�b��ŊSp�l�Lw�ĂQ?�Mȳ����}Ig�a}C�!y��9��ȯ`��ן\z�n�ϥL��;-��k,b���׈"-k)�u�����hq���0�tk��%Y�]�sxa�>�I�.�O�9�cU����HC$ߪ�&��	b���J��|D�A�}����T��Q�Q��	䢃Er~����>�'��$�vq��
5E;!����cPU[p�����<�AsRu֛ZB:�W�J�`��g��\ۤ�)�dV���7gZ	�F��j�,�TO!p���+� 򳊅�<���C<���77�A։�b���}�S��B�a`���/���Y�C?<�M�9Q�����{G!1q�[��J���@��!*]��vF;B�xM�%<�̸�v<(q��鮋%�����9M,�z �cBFV4���ss|���#�>%���&�Ad$a�Ϥ�X��Z�(���&dg�U�;C��M�p�@\9�5V>�LӴ��
���J�O4H)l��:_�]��N�DV�>��h1��`�L�2<��x���\��ܹ"d��2s��t�T��4ߢ�|q?ȣǟ�%� �!��q�Q+���lz�ǹ ��S���:<�!��`��g��g����-t�		/]�@� �ZJ�(��qx�r�A*@KW���}߮s@���A��k�Ȭ6��ZB���r�o:�7�~ƙ�N�GkTָ�-�[�e�{������p�%rt���5��/��?�@:��GRZy{�'�Ht� �bbs�]�V���,��Ÿ`�7.���S�o�p�8����mFMa�v���Z~�26y��B�"3�V���}�Cv܉ߍ����/��\����X�X擖{GU�p��bU� y��l4l��jaߧ�Z���r��F�|�^��=�&X�|�
�h���;�]p6�)�>�c�s���_/� `qXy=ih{�~��|�H��/lQ��mf9^m�>�C#1a�B���_O�7�8��$������h1��u�I�RGbB�[zB�L���I�k��m�#`턒V�a�SYsP?��!�1�q�K����-X�oDa$C	�P{�����\*֘e�J�Z��������R��70>��K�����(½p�����H_%�V��*�k�i���8���3r xH�ꔎ���e��G�SΐI���/�E�EG�����0b͵M�:mN=��F��qXf�������Vqw�lY7��{0Hu՟Z(�r�"61k�y���՚E��j��rp�b =���Zpd���?}?���}�ŝ~�� �vj��,&�s�!��V�3:��/�]�7,����*�����' $8�H��$d��5O�����������B~��D�N�l9Ե���@�G�Ֆc��y�>`��;"��p!�i��WW����[9�1�z�ʳqe��R���˴�Z-�Ŷ�o�̭�X��D;����lhqx�?2áX��7m:�чҒ&ߵ�ۂ>�����9A^��a���8�7;Z��Y�fc0E�����a�@��E��٧�x�&"�l�P�)D��
�	�ϡ�]j�� ��<zm��&R��!��H���� O?��͗���*b�%���?�`��<��*[�T�c�����c7�|W_*F"񪄾�@�ym�p������ J'���)Rׁ�@}sB.e�ٱ�ϥ�n�v�,{a߱�Bf��~%��0>c��SN�v���IdH��í�G_؆gn"�f�)���;�m�Ұ��������Ŗ�M���0����).݆ҋ�HJG��x�s.� �
�&��j�&����vu�h�I�����N��)�Hrp¤��j�씹X��OB�3_��C`��G���QW�R������Ky�L�Y�Lڒd
f��yґ�m��YKd&���S�-1c�°3�q���?el����5 �d�}����0��'����qP�҇�i��nxH�f��b|�aJ��#s�Je�c��L�a�C�݃�~�n�?�N���D&`��,��/�S.��w�m�2���/xO��0�3�E��p�K8"V�A2p�j|�ykU��jg���f�h�m����:�nd��φFg��,�1@t��	���a����ҥr#�@f�Ȟ̲3��
�Jyդ7y�M�mgA��t،�>����	:P��gO� @ۧ�><�&�x��/&)a�ja�3�ع%�1!����ڗ��泂��B�"�P�M��C�0:�ʮ
����C+
ڕ� ۃk
��6r��#D}���(������@�a6���P������[=�A��I��M�
�6בZ.s?��I�J����3c����M� ]���q�M/. �R�|	��vѶu���@q��\)^t���ق)�k7�
R�(�?6���y���3#^�!����ӷ��9#SS_r���Z$z'ْ�-�i'&�0򞺷��,%ʬ���_��}������ָ䔧���V�m��,��l�Pj�P~��� 7)I�f́���iHҕ�ƒ���\�+�H�f�7/�:'�+fp��qi�� pb��j�o~���1�����&��@KQ�{�ɚv��}g���Χ��Y�������r7с�4�����7.�8���}�6�>��(pfTb��4�@NH^������V�Cq�@3x�3� �ac@�>�w��WF&�TΈb��ON.Pe���g�1�`(�f���wU��`�5D:=�4���� �)��~TN���@K_��V�ӷ�Q��-���v���醹�38�a#�깝�����L���C��#�&J�~����1j�b�kX��;u����1Y���U��jwB��в8~��(�Ml1Q$4��z�
��Pe�t%TG�n�x���O�j���%�kM���{Ai
�'�iI0e1��:ؤ
����fԛJ熎��w�s���3<w疑���_.qu���h�y���j�\�b
F�P9�܊�xo��cW[���)UX̞(�V-Ɨ�
�w�$	�����U!rv<1P�G��̱TŦ,��H5�\uL�Knb��u���`�B�C�B�YR��Lda,�����ήj���|w�5�?6�X�"��e�c����o�6y$��p������h��e� +E��r��×����	*��5 �]y8_�>,kIc��yͮ��r��3[�OxԄn��c���i�!DJ����x7�8@�We�	e�o ��D�p�+k��<��o�ue=^�z��������yݩ(���ߴ� ��S�6�3++(ş���$W��06z�<iJ�9M��}����l��v�� -�\<�mFı�i�����0~�o���d��ߵ��̅w �2e��.!p���+f��1����2�
��ܨkug���̲dU�\@2�ۮ-5i����� ���]] \MDCl�J�n�Ed4�5� ��?hs%o�(�^[d�����(��&;�ZZ�=�R��qF�4A+.i���dfW����c�΅�z��$��.�N�v�Sҙ�M���� SV�^�5�9'�軡��A�1�O�2�o�����4r]�܇q���u�(EmKƀ%0�Q��J�9�V�;Wd��{�'��3�?���l�ȁϜ(�Qy[��ǚ��Ɍ咩���$���:
��Z�\�M�2��p��Kl2�p�cF͚Í���a�]����J+�ilO<�G� �#HZ��W�\	���Lo8�۟�DTσ���F$�Ov�_�Ԓ�'���&%��c3�
�
��8��>��u�����x��.վN�����n^�ҷRcu���V\���b�2���Z�e��W9>i�o���G���z92�
��W��m���Q���	#?���S���j��$v#��Դ6:z��S�>ۭ�ݴo�L�KjH�p��.}��x"�ح�w��lP(�Q�ɸ�phe��Ѳ�K�}�9�
�׽�'��:���W��?\��y_ A��_��a�&����Ꞗ��Z�%P�S����zQ��@s����nL�����ż�🉶�<�;�zG�R�1�p3��&r���`���&��?ى�sz���4�z�O9K�;q:盺�E�����Py���'��z��_���� �G��}ŏ5�
�� �RC
ʺ+Ϝh@���E�V��F"�K�t���`G�60i��9G�c ��S
uL\� �<Cڅ�������lt��sYL��4q@���X�G�`*j�<�\l��J�oT��1�T�
[ f��_��Ƴ�
�3�F���H��;��w���6����Q�O���/��/T���3��p7�4v��YC~�.�]�`L�����U0��H�_�lU����E�C�!,y�0HU�@���{m�m��to�ؑ�fS0��?w,���=�����i�=-���<�)v:��b��$�����Q�Kt��[��{)�!��J�"����3����r��3�B{ijҐo�d�E"j���?�{�)�3����Nk� ^�ǀ�*��_�����ϊ�y�g��F)�5����t�ڨU,�jŰ���蝏yb�BJ6N�@��&��n	�$��0�9B|��I�..����K����Q���CP0͹�U��6Ŗ��Fc��%����TFa�	�_�ErJ��rWX��H����c�7�/]Y"�)~
��N�[N\L"y��p|���4�/H�L����#6j�*lD�^��Ehst��G��{sEJƇ6����ͼ99��|�gT���c�]̊f1N���*g\4qv��IЊه_�/MX�F;��Ո&	p��Q>�	��!��I�3�f��Z�Z��)H����:A0o!hf��A�t��M�T���VW��ɯ�*�^R���b����͉l'~LC�(2��`�F��C�%����o��sR�@͏��3" �5(e����3��ekdҥwY��S�,(���ۖ'Đa`>�Y2�H����Ɓ�!�c	���>�����$1&��kt��L��c�opy�⩮,������'��l�|�9K����al��c6�~�����H��/�a0��2M��/s�.��@��TǹF�4`:�z�&"K4n�96�Q�Z9����(.�)#UM�`��{׹l#rSV���1����~|���.��<�Z7	�+��1_V�!�~�R*6�=����czS:'���=�)&�o$3�$n���+��I9��n��S�" h��/�L�j)~;�E<b)��|}�-bWx����.��ƨ�ԁ`����O�ߣ��b�eۥ����z��-�R�n�@��J�`L>G��݋�,�T��QGAR' [�ӽ��<�|�~2����q?�|�uf͔���	ڗ���C$ �O�����*t.�b.ߞ���?"U�7�J�O&љ�g��������+��l��.�,�ϋ�-���ND�l���O�ˬ��4��H�vw9|7آcՍ�`ɯ�Q���5`�rm��{�&���#innv�xK���[C�7����y��r ����Z�ߑ�J��ʡ�L�ߞ���9�p��C����R���G�;�M�* �H�	{i��^��F�#�7.�=jR>W���*(<��yz;����(����ͦ��O�=9�k��!����+%�P{!D���ƪ�����/ڠ��D�)��Z�$r��{1�9�E=}<�x��p�!zj�n�0p�A<��,"Y�3�����'tzmM��h��}�HY���\�֘�fyӑO�8_�H�ݽs�:n�g��E�^����4�+��Az�u�L��*^�ؔ����<9�Ռ��W
�j���b#J�t5��M���T�����B�m�a거�ϥ����~.{�9�Y�z�����3�����3%<�-�74�w몙�Ki�
(!e��?���9S��ލUœ�C�Hu����-ߣ��t;����),�w���P�n��n��Na�g(wf���5��0�N�y@��Y|�7ز���_&
�g����4\@0i������d57q��>�N.*A�^��P@����r	ݝ�֩v	^K������{Ԣ�G6V��y��Ds��N��˴O�ऱ�>FH�+i���8��6��$�-#,�nm��V���N���D��ko�K�@Li���.�E�mS�q<�2� �����bVS��1�1��b��>4W������ð>V[z�������Ǎo$��_��yZ�e��\�Q���X��U��[Eo_�$�b�AI�T�3��s�Q�Fw_<�JШ�#�LM�w�u���G�z<sa�ӗ9z��� 1H�X��������n���c�~k��~7}��Mx�8��p6�_�w|K>
�!�5��#>߼�E"T�w�7���֯���	��|����:!����>�m�+�+�%�A���#���6�2�>'1,��%BZ˅��5�(	%%��hBژ�.r526.I��WH�E>)��Q����M'�t��s�_ȼ.G�!+��P��Ll�6ũ��L�f΁��렑>��	��ܸȰ�h�{�ɖ��4È�?M�J�ʥ����zsv�J<�s�Kxb�ox�_�qL��	8p:�:N���)�I��e�Ď� k���wش���Ň������Cvd�@��7��:��3N�ȓAF]X҃̂:6�-��`	b���_0S��E�zɻ�{C{:C��a�>|�]�$�Q�Hq��&C����jfSi�����!w�͠U�����G 0����\�����2�<ru|6`��)�PH����7��h���o:�P����bZ�e�Zz?�Ǐ*�$ρ�ܑ�]������'b�LJ��$���a��]�M�Qs���u�f�T��A��F��9�$�HUov�`Ec��X���?��-?�a�f�)E�����
�WT��}��HѪ�.��4��d��}��d|Zh����
̝�w��M
#t�BIC�#�d8|/Ѩ��K�^��#|����K����7&��I��t����0�V�D8A��M`��S��uɖR��ӟ��c����(�wq.j���N�狂�#���z �;�XQF�W1B3����/��ػ����'����mtuET">%i��x#�C��R�6o!��������o!f�!�A]ꮇ�5�c���2r��٥�w�5>?����ALveq�h��\�6nH�>������s�4��O\��� 2�k����|i2���j��Sq�&���y��ю��̤CV�K/0;�Y�{@�R�x9�Q5֝��׷.'�#����*{����
�b>K{_���xc�����2$;A�]�s��$�<	��"lc�^���$�Z�g��3�v`�Q��ZGX���KE�^�HN�G��ivM*�e?�k�޿3�'5u���ܔk����ֵ��`* �]���W��F(�Z⋊�7�ܑ��W � p���re�����4��ڱ�An]�]0�j�KBE?
k��ۇmx�5��uS��#��-�g�!#@���|��j1�x�*
n���b	n����
�h������c��/��N�&�x����\4�z�AX�us�|�=�����)nł��Z�Z��A����P#�&�w��)�m�! ���0���>�t�rBL�)���r�<&"1%U�s(&���?�sg�0�-_�f�l`���$K�
y'��<3G�e��Cɉ���r��V$[�>>U�a��ds����:��� eXt7�T�R�����\4�k�Ѷ���-5�8ov��I��D����chU���'�s��j����,~�;��QA��I���n� uo�l�u�4±�ْÒ;'cz&-<�1�XسT�]_Z"�G?C�|ʪ"EASO��5�QW���AG2���f��i���G����?l���ⷡz�����H��^^(�JpH�֦�P��7�m?=^���18=������=�)�yd�U�4?M�<g;��秏��c=N7�4�p�ޕXe�sZ`٣��Uj�=""k��%Y���z����?����欨�'��}��/g���md�q{[�hL�w���K/ϳگ>:_3{�F�0G�[���T�Pi=�C5ގ�i�#e��©JT=qg��Iz.��L��	��z�1?�־O�q�-�c��o�G0��8��<�v�m������ �7�����{wc��h�Hg˝��+ѱ�b냄tYz��l2�W
��*�����B�T]6+!l&�/Hw��;�,�����Ƒb[Bq-b���i�p��EXJƴ �hͣ){Dd<x�6O�3(27f=��<�����'�ZФ%&0��B3��'8�hO��p��KVe�՚�C'^�@�z�◞����+7呢=U��J�i�Ŋ�iS��kPd�=,�t�n5)\�N�) k+\=�&�|��U��p����p����&��[t��@7)��8 �s�EYB�B���A��t&ha��<�a�=�>*�.Td��'b����U�P��Ƒ��$n�~~�I��u�$�{��{���f�3\�X�1@s�_��1�B��R���?ݴ^|h������(��3�P��[a(�d]�L>�T������{�C;�,N�(�q^�� 0���
�"����Ǽ�(�;6F�R�}�T�Z\xW|W[8��M�n�e+���fP}� @�I�l��� �}ը��=�pG*��Z:���oѵVIJ��=���|�{�z��w�E��nE�_���^�h���������'�O�RWxx���=���e���C�Ŏ���ą�E�QG����Wp��	=	j>�����5������SmoAS��1z|��%�2aW�+��2`P�>�e;�D4��Q��5��TS�j��[������ˀ�:Z�p�f4e�#W>Эe�ڨa�h�"�Y4��EfّF�ΣW�����������'�3_��Ci�p�Rx�q�B��ɚ3ښMp-��cÓ!�\�D���y��ɒK�Ej:c�>���&Bp��[��A�t��d�nBxX��~��f�=*� ��2m�/�B!�M����\�)�[\q�5��$8�l���)�7����	,꣚E���0���-�`����_W*.�E�������C1S�=�$�5�����չ����� h�g�ȍ^���$�F�u>Si�ԍb?ҍ��VX��)W�3���۵`����������9E�La/�"n8Fau���K��!���3rĶ:�� ��5��s5��ǏuI2���9<��J�B���/AId�W�[���v>!x��B�lJB��l>�n�������7^�Z�W/]�M���))].����Ξ�:�c���@S�7ʖm�\��C�� N���\��@�H��ݪÄ0�i��o�m���İ/R�ܨ��$��6�_�>h$����*�;ܻP+�J�� w��}���*�.��d�$��JU1@���i�n�Ad�^��n�����%y�|8#�6�� }��U*^u�(��׼�X�k�'��>I�j.�w�����=��}���g�/Z�f��B=�F�4���UeXN�E<61V�G��>Ԙ��/�����d��p��y�SGۍ�PT��k6�{�Ÿ�ū���r[{Ϡ�MUEv��j�E	����q�Ir�5c�Ff=�h~H6Au9xPԥRS!����ω�`����/�0ǫv�x��PDU
�z�e�`��5q�p��[�y#����F7���Gf������7{��?�H౶�"�ʔLP�w�
�R�L���u����MR+������O�	�N�F�f����:4�_[d~4j�hI�J/��#�-�k�Z�ʸ�Y�L,�Ϛ��%���qĐ`�ފ�f��Zg�|+��ZsO��r�����0E�����cy<BC"�˄џᖛD�PO
�q�Yf]�j��t}Pfj�S��Nc%��>f�)|�!�ƒ��]S����!�C�7��u"�Q9�:��=�E�+�?cRL��ի�A�'���:��g�wǺ��C,�3�,AՔ�d���6?�3�E�U���4�vT��`�����HD�w�N�X1	�� e��#13.��t�.ν�`�p
֞�uE(�!P����Ъѵm�q�*��~v�6��e����J5q�uL�g����X���a=�d�O��1�1����>3��w�c'R���Oe:�aW3���ʬwo呰j�q���?����B��4`Ú ��Ћ0�X�K�0��G'4��1K�u�'�x��Oԟ����O��e��g��}{�fn���?�����,�.��P��_W@uR/m=u�d �W��`_�,��`0�G�,�^�E$:�n6�!����V*���MS��i!��dw�ؔ�f);���e:V�I��(�r��)��KZJ�˳�+��;yR?���D��YLŸ ��RS�	�d����|ڜ�#��W���@,ן�&,�^�R�gA�XU7TDcK��WkzzF�}�<�2��*9��
o�O;G\;�R" ɞ�uf�����lသ���_V&&5�K1GO�x�[��0"�<����Ĭ'���~,�u3Z��f{�jڠ�����?��w�?�W��@b����ů���^����W�<f�}*s2�?��IB��G2�1�����~�6�O>b��A�����5�}~ fdp���Lz��|�"E�=���Cn��]��0�'T�m��=�t�t�
sv/�E�XD�q&��r��'�;�v����Hz(�������S��u$F�9R����Nl�~�!r�b�k�4��L�h�^^�Wf�z�����2��x�wI!?=�#:��@�ؙ�9��P�6@'��A������*" %����z7d�
?�@��C���Q<<�D����,K|֩�d��d}+ek��a)h�@07���GDU�N�/k��KQ��(�CD�l�r&0�*LeR�T��8�)���V�������Z��㢃} �eTE�9!�M�Ȅeȏ�|�W�뒐�O���GG��

����6^�Fo�~�n�$��(G^C��x�̾"�W�l�t��[8�ul�C�
�%���I,g˭$ /�?J�����Ia���� ��޽�Os�ўoZ ���hw�$��;e�yt��/�Զ�NߏqU��D��+�a1	��� ���`D(��|�'��+� G�Τ�ߎs�z�7��tG˴�)�4�I��@��#g⦢
����r���p�P{e��cӣ�͔�'���Ԕ�A6���Y�p��K,��۩�y����O�1��s���'��?�߽�.d��PgY7
>�س%H��X� J?Z�ظ�	���E]>���%������LAN��l���Z��z�,�{�������
��+J��e�����m������>�Vt.�Oc-���T�K�.GĈ���+;�j�C��w�$\�Mcl��9������X>� 1��q�݋w?8B[X�����_ʹ;��g  .^M���E��6�<��Dm���\b7�,ǉ��>1�;��ie�kÉ�ur���gI�joS�f�U}?q{8T�r}n�*@ַ�:ɓ� �"0�%�;�� �����YZ�u�>�ɭ�l����[����G�G��tQ�>q=eЉ쒪��j(�<���_^���0c�ȇH"dy{��8e
�m&0v�M ���p��+^����r���Ӏ��Jy����������:�7v^F���;S�e?G,�>U}/���-ŧM��X%�l�Z�-(��2��X��}0��Y���G�	���(J[�H�,<���l��v��+'��*���I���;N�s��&>�1�u��H�j�d�mK�+banA�-ųdů�oƯ���,ʒ ���N����	�o�Rϋp��(X,��ޓ��|iM�'n�O?��_	Y�}�t��BdȔ�	����O;��MD��x~[�Wҥ<�TY�T�䊫>�1�Qd`��@Dj_k�_Ǥ�MW����>#���7��$��5�C�e�\��O��-�����:�5�����ـ,�s�� F5�D��+)zIG����L��*��B����8��y���IJ��Q�L=e5E@�&�G���a��ZJ�Ul�+w�*���g!f��
�b}<7�<�%�id�J�	�!�\NT
���\[��]q��իWC����]����]3/Ի݃�m�=Kb�9q@&5�oYN�Of�O���O>��>�m��q��S1�6菂\�ș~:���B]do�{����E�������y�����K8#����̫�P�:��;����GL���b������V� Y�a��^\�o�+Y� ��^#p#L� �H��?nG��� 	�q���.��y�R��e]���� �m 8���y�R���e��7k}��`�Dے��t���O$1�o}u�L'k��|�9z�yg�ش��:~I�r�[+���ť��IY� ��ދ�_�4�3�3@���Zt�>�VX�- �]f�N���Ls���xL��=���py���:���\������XR���
!Lʠ!�x�5qP[U�d3�z<Sե;�Ceq��=Јܥ��q���+;O�N�Q�l�f���i���ǿ��J��C��j��b�#%��tO׾�������>9n��&>���j=߱��^��8�����=�T0S�aO��g�jr`�[�FM��FA<�%!+��^r$����Xu�cܘ����q��
�~77�9>!�11A;ր�A�B�Bo�#X,%f�[WJ8pX���n@L�,��~�KA��:����O6f�h+�T�f�����̵�l8H��%nPz8.���]I}��������Z#�#��-m�h��8':�1��w�V����A��BPY�rI���A�b��f>z%%��$zzR�E�Z�~�И�&PZw>�?D��Q��X���M����������cH�4	V�H�%����I 8�C��<����A��Oc�3X5?�ZXC�Qw	�n��W���zU�1ꋢ4V�Չ���ytG@i�Yt=�Mn:��?����aP�A(�
L���d�N������^g}�i%���-fd�?�������?�	�u�1,����ce��Z_\n�
_M�����w����ͻ���@lS�8��Wb�{'��Co&��>�
�2�"������C���=�K#������� �J����e�y�0|�wgU'�6�( <�j�R6/J�Izf��ٔ��Bc�����5-s8%��OW<s���ݲ��\�{�7�Yי�q���wY�*�
~ؗ�ն�3Y;2'�	��6a�s�B��s�T��yI*�O;/���?��a3�Nw��L��#f���
k�◧C�b���.�g���!����~ �����^ ������6z��!a�E�qWۭp��1{�N6�d��a�}�k�´~�/�����&�6����gmeZ^�����VqQ��E�e��P��e�.q7w$�$�K�Yt�I�Ry*�M[���+c�m��!+z "�Fn�������Њ���@�9�(��X	ƹgS4�H����L\���*�iھv��֡��$�b��-z˯�,?�ϲ}9@���g�V�<sw��ġD�s"�J���ؖ�����z*KXh��ڙVɠ�o��z��z�V���Z���� ��~�O2OJ���U�/�֩� V�n��v h�F<i�� �Z\�@ʛ�.!�[.��u8+�1a�W�C���>�w#K��������i����>E�*�XQ
�Zˎ��&�lu����[�Js�UZ�3#c��Fo��cd#�����a����sS_���r�
WQ�fw�+|9-�D�0��m�t�����ZtT�]�Ha���+��u��,>:<r�&�XRʢ=�oGƄ�GϤ�WU{�K�#ױ�cX.|v���U���ICԗ����Rʊ#�Q��i���������R�����Ha��(��;��lꢺ#W%Q�ΰ�$�*��Dwhw���t�6��Cj��	��wd~��v�F�!��*w���� ��CC�uJ�5�9Z6Ur�]�FIXϳ5X팰M%�p�,�S�ؤw""o�,�;�E1�~������d1�/��;hs����hmR����-�Jۙϥ�]{�C���إ��{��eg�W�T��L-��;��݂�3m�j^���R1*y!Ѽ��
c�	���{�?�T7lE|L{K"�wؒb�
"덈�`��5�c�yu<��z�{��/�ϋ�e�=���v#/l�����|0vi�-2�?����$�OƠ��6-S���Mqb���kB����Gh��S�'֓�~���:��R�T�D���l�뱈p��+���wS���r���3�s�c��z����b���Ohs���>Y�䟒�y�.���(�2@#l�J��I�����:1)�{�!���F�Ѐ�OxQ��p	I$S��N�;�#����OR���q�|���(�)2�����\�|��o�G�=�Ag8�+޴f~@��D��4Æ�Va����?"�Q0���}��]�� ����z9��9���A�:m!r�iF0ߗ��$�0��h�Bʝ�̸�Xɱo�ﺵ ��VF�0�}���m�$�G��;@t�+V�ռ@G��)ƀ8ؗa��ֲ���F1H��*�u��U�������1.ͷ��N��*� ��3��\��m0[�E)*�U����O�=�Yn	K�eI8�SLQK֔�����m�TY�ͦM��0�zg+��B��p$�k�Ͽ��!@Wݨ(@��^QL��=��m���%TI)sd�NO ��pX�fE�K����V�3�g+���@�r�����n�6��ܪ-K�b����n�?$���n�Le#+K�h���ч�54!Jpkr<�������J�1�ˬ�+��9�`�{U�ˁ��-.�z�L�Mqm���P�C)�����f��T��*��}��r����3��H���X��;~�����b��N�1����6[X;k�w��d���|��Ȏ&��D�N��� �n)J!D�����7����QT1�y�A�CU��/п7��k^{9��О=� ���j��pY�����l�ۘǕ��Q'-W�����g_�[�$~���#�Ԭ���\��ZI8C���aG�)�8��эz�O�B��A�^]"��,+3e�<ㆰHmb��M�\g�E�8~$9$��e�<l�5���@9�9�~�����;L����38�F3���:~�35�������Ts�j����|�?�9�D7�/�������Գ�G���3ZE-K°�\!���!�(���
�n8�v)"�b(���#�F4Sl��Y�!��S�eЭ�C}�/��:�dF����.��]���<	���9��֤��-J
�-�\E���U���\�&b���M�|�_���9��,�|�k�t�1����ْ�l�<���[Ym���X�+!�r��:�qb<H��rXJ����VĿ�����]#��n�4UZ� �8��$����cwf��;��~g�^f �`
J&��m�5��N�		���^�0�:��Xxf呬�Ir ��O}ĳ �&*<^3k>��]�騝�,�ǝ�jg�i{釮j���Z,O��2��E�[�CK�v�]eK���C�R�DRS7������j�LS�!���X��	j�.�
Vz��BK�^_��9ς�"��#����:��g��a��3��(oB�E_Ҭ�g%�=zeA�\���p�W��WT=Y�A[�t��M��L�ġ�%���Fa�]�x��}{�����N���5�"m��ُ�_��;ݝ���hd�,h¹�Ɇ]$���/�cÔ�=��#�=c�L��cq�]�c��XX����=�BIS��=�D"��%�uJ}5x;�=������?FǩZ��&�7c&&%�'�P4����i*�P�P_.��%d�R����"�笤���	сž���1���C��o����R�T{rW�u��]b�vB
�$�xah]�Ͷ�$��20?�q()��������õ��Y{d0,�V6�� ���Y~N����x�H/Į��js��b���o!�b6�Y<A��� ��OXRI�Ɇ��'����ojT���z����',��h��2��v��qV\]���N�%�ZMONV`�	? X#G�3������Ra��Ѩkl��8̪��0S{�d�%R �]���J����܃[�ʡO�K�r[�x"����7Eي�#8j3i�_��W,�D����ַ	MZf���T�#���ݍ�i��!�e�X�)Kw֔ʺ-�̍���P�}Ii�(��B�B�rY���&s�R�lA�Ď��;t)cц�H�	IftWK�a��jrVl�0b����	u��B���T�G����C{Uc����/G-s|�s�=u��V��q��]g�:~��[�u|�:W;2(��m�D��\��&A�,��p�UGS��K>l�*	M�U��AC���,�7���XCf[�F{�y�V��ϗ���@J]k�ڧ6��OS2!���C.V�h�8/?B�%utF�'C�~����.S��&8�E_* Z��XxF8�V?���n�h/Y�P �s�f��`s��`7;�E�]�m��@�����=�	g���25��fZ����UiM�m����9BЂK.SOc���m�DBr~���O���$��k��si��_��r�dtBm��.��r1�qН�+]"#�����`Bg�70��tBb���_�=!��]�MSY@���a��u�}a�&H���NW��'߈b?��vC��|b YdN%��(�
7��!�l��
x=)0�E�$������<a�B��z%S��_lMh�u9�H������޸��u������{%˦�x�ǎ��1g�e��W�6{���n
����1�����'�A�WF��<f6�k}�13�F�%�5��IVob�4ޗ,B.uq
ٗ!��˔DG�KU�飱<N�P��a2���%�tʟ7��3�	�-�7��� w?M0�Z�y�E%��˦�5��Φgj��˄����}�[c�E�����j"K��&�ʣ���(IЋIB��)�8!#l3��T�vtN��X�p�������:S�N���A�c�u��>��v}ޜ����e��^�l"���C���W����@�蓡�+5}�����2�r{�7>����U{i��b{�bզ0|���q��9Z�E�_�G)0~+�]�,�З�7r�5�Ȱ�2���,-z�vh��+Dl�W�aM�/�����D��ƮŔ�)C5���a!�����0�����,��=�:T�Z�$`%���_��7�(p���Î����&=�-�n{������|&�D��E��J�:Y�V{��k�ZH�O�CmUƹu�:%�D+�=���2no{	�z�m�}��IZ�À����y*S��b�����47��Qcɋ2)0��s��Ӝ��Bs��ܰ�=�&|�*���f��JM��/л�qT;�'�nӃj�"���:@i���mQކ�@8�[W�Ϙ%�0ne]��˦ҹ��D��V���&�,Du��trDI>�B��EZ�>~�X������O�I�Ģ����E�rǡ�˷�]�3F#�v��P���`��@�K�Q(ﳈ�dIjF�Q�`ֈ�Bŵj����r�C{+�o�r�J��:0�3�*����ʔ�q�d�:�k��%m��4p�B^���ign��a&BH�bS�:4G��Ӕ�ɯ��B(�}�ly��*����|q_e&����1Ew��'φ��`��rq�����ګD!�{(�ٹ��x+S�o@j�Ip]�� n*���	��|�B������-�i2#�*�FXP�<hy��wO���8��޵��W�X�߇��~UK�X{6\�7�l�"L�n���y����� �~���ו͞i������'��f�X��J��� ��&D}J�J5�&^��l ���+���6��*k�Af�W���1�����Ԃ��E�$:��8�������}/�Q����q�V����N����1M�"{c���X�3����x��6�O 90�щ%�'�A�7$�:��d�l������2�qZMn�
he�;ʯ]�z����2��a��x�ҵX� ���ئr�{^��V=ٓ�h	�X�g�,�֑�f9\Ήɔ>��7Dc/��сfk~[!,�U'q�H?-R�oX���d�����s0���
 N�`��T�O��-��8#�o"C��m(��v/���ȭ���PS��	aV֤x��
�Vyh��r?�w��pn]�(X�ף�W�(g����� H��wꚷ�� .�[���e��s_�^C����s���-��7���
�r8f
�`�qp7����:._V������{j�[tثa��5;� ��<�#^�_�a��J�o�:��ָ��
y�=^Ը`u�A8��,`�1+s/���V���u
��V$��Y���q����&gs�%��gt+���R��gg05���V�b��:��J-�I�&;C��i��k�s��	L^���E��B�)����o-�X�8A��*���,���
r�B�ڕMĴ�F����\d ��6j��Y6�ۺ��dn��"=U�r� ��K���N���A�D��!�π*�Cqx���pټ��������bN�z�:�],�>�(��{��EǠ�7�1��T�p���RV�C,�x�w��ы�����R��N5�oŃ�X��o�� 6�^(*��v�DUg��#��;r��� ���9���𰞤X�2q��2���u�DE��X�*0��nk�N�+����s+�17�Ԫ]7B�;#��}NrÓ.7��-����O%�q�v�^Hu��o��,ݩ����i�A�Rq��2BXʼ�p`)#��Oۚ�S|��ZJ����?�y� �����Jo���H��rn�}���(.;�!�LX*	�A�I�{�pj
/�q=$)�5���l���x��Z���*,(4��%/��TR �/�LC�"�覃S�Ls~���%)+=5��R��1eΓ�S��ҵ$�~,��Z�&��t�~��w����d�������ӝ��`�l��%Q$�$!/��{Z�!����ܠ�v�&�<����pR\-_Ն�|�h�o�5hsn,�����w�5Q�A|�j����|�mru����
��\Q�v�ϒ4�v��~�9u�l�� 	X�ޟ����m���ԇ�v7K e��7���h!�_os�7�#�[V��\��b&��'�@_$�����Ӓ#�+>�����
�=�_��^��|@��Lژ��X�D\�Ȥ�2��bx�5d�܉����ś�P�*�MF��e���&�G�}}�6��� �ے<h��nz\}7�v(a}D�`?)>�C@ �ܨ䟔��;V���.)B�A��*���2z~l�OK���&�U̡�����-لY(�p�GLÚ�_�q�e</Ԫa��ߣʋ�S��}� R�����L�42 ���hI;�N�����xn����<�_|�tD�u�s��@Z�`�r.�^$cN*��4����Fm	4�	fG��rz`؁g��@����U@))D�߻��>D�Py�W�SO'n�,mM2!�;��>�"����0o�N��$ۦ����K$Cb���f��T��ͼ&��y�\�괺�����+=�F׭a��Ee���=xW0�s�̔
��ß����HBV�F9$̛�`�%M�h�x�|�%oɭ(�������/��Ⱥ[��}<Z��׃g�X���UW�OpX��,�|OTt�����9�-z�9Y1�������z9IIv��w��$��qgx�+�mww���љҭ���:�y��Z��4��x`;����/
���͈���Pݵx�:�ֿ����2dN�]	Ǉ���YuC��d�&g4ʈq�s�Fw]��ڟ��Um��T��H���c>����A���p\=G�y�so�#{�O�m��\;������τ�g\�aO|6�D�z����.	�Q�o`��),�F�K��o�?D�ֻ�\6:��\5��}�B6�10y܄�a�9��>��ݙQ�T�WZ�HwI�  I�H6Єp���ٗm-�gIЈ��Oq��c��� �b������xa䯀��+eC��L7%��t���a�Ǒ�$���)h#�����#�|��!TdMb0k���"���õ�8[;M?5�����g� �>�<!Z�Ֆ	T	���[�Xx���R"�%�N��.~`j�k����?�Kp�M�x<2���2�8B̝G�/}��rJ�Ƃz��nNFo�G5��S%���ل1���$��ĥK[��)��}��*�O���!�i���V�L�~IШ�g�e�+qA����8p�րd��IQ����ʓ݂@�-����Tߔ��nU������z1P�r�X'3GV����8���-�&h�h;t�b1�.�J�K�D�ѳ��ʲ�Ӹ�>���CC�ʃ)���`�`���rkq ���f�.[Փr��4�v�\��!v��a�u�D솬.2����M�6Z�L��J3�m��;������ꝶ�|�?^/4�5��A��#������c`n��1찍��
����A���34��?
b�M�P�	� R�#��	����O��&�tIP`��jn	T�pQp�'�ە~F<	f�.];�Vp*��Y"��T%�7R�Ӟ����KF�_�1�,�u�S��r�C���qn1��ݙ�u�~9��֛c�Y�g�#@lC�a�y�}�`[����\�G��Z)3���?�`�����G�>i�U^�ڞi��;և���h�8|���P��}��ִRWyƸ�Fi��J��}d���8�4�z'jC\�jp��'�"�� ��O�����!�-��ÚuѹgM�<�ڃϣ ��srդ*��zu�܅5=��dbհ+o����;�	Ok*v����|��$'�{}�3���m�x^C�}��eM�#߻�	z�E	:��U��G[~+@�H��*���j����'P3���Xa�g�Ǫ�a����S<�@���qٺ�-�Qӳ�_�e�U'�����k<�{�v��4���浑�L�~)}gQ����X��7��i�D;b@��G��@����� �̹�B_`U�e���x��Ot�	��Ǭ��'u�i��3ߕ��8#�55N�꣭�cI؊��d~:�͹G��gV��
��搌h����=�=�u7�'�Q�/`$�H�u|e4���ЦD��ucp[`���'��»y�����=O4!K�g����5 )7�'#m`��E/�W~�� �P��ו�k�'l��}n��j�G�R\�0|��kLlFU�=���[�w�31Lf�}\�	Fc�BC?N��5��H�T7��R��:V��3C��$��`�K���řZ�~�.���m�Q8�R�DdT��z���nH���gN�ܦ�P6:>�A��G���?�%�?��֩D,�}��*���x��Zc����g�^��K��		{z�eJ�?��Y���s�#f�	�#�Đ�(.��r/&����i2ԆfU�;�v	�%F�5�_f�g�Ny�D�;�ý��nu�+)��U���CV����:�Q�x��ܩ;)m����K�$��\ܔ�7W���
����,V?�=��8�w�DFyZ\4A�!9�)�@`Wct�d�1Mm~]���^qu�wr kT�/�������}G2p���I�qddm����;YX;��i����2P��[~��9;��ķ@�б,Y*��%>��󽝤��^��LBi��
�ck[��ͥ�Nz�?D�TC-Զ�F��������*�	�ꁟ��~J���뤌���R)�����ɧo�� z(Ų1�fG��12F4�p��(���{
+���]���W_���D�@AʡLRY�C�c/�R}念�{]�g�^�i���^mfD�G�������
��d}7X!�݃R,_�+]&�������w��bx��Vy��ӋB�!���	�Tl B�&])��W�j&O}��Pu��:����
�<��z�dxz�V��"	͜��k�´��nbbV�w�;����H�����Y<�?|c��F�S]�� ��E�RBΗ�V��%F�x>�8MA��/�N
JlAx�H`��z��+i;7�<;)��+�[>Mglu�@��{��.��'�A��P�q��%B�#��(D RoR���?̘��P�9�\�~�f����8��چ�-q��hd���gD̝ɺ��������4���;���(��*FJ�|V`-�O��\N�z�qs�׈-)@[�*�NDE���?P�P��O�y8�c�*��:8v��[�-�্t�k���BN'),Dػ
�h~xI��i�72��A�,���P��N�*�3�bŜtWQC�����(8�)Dd�乎���AK�u�ӭu��f����>����ֆ���LΔr0�*b�]Ńy@.<��Q\���ˠ��vkDꌄ��\1�� Q�������v���&�`��F,f�,[h)1��l�ǬO��0��~��r91�j�*p� Fh~��/c�ڜLOa�r�f����߬}���	$�´ň
�.��W��N��s��N�
y�q`�S���6c=�+b@.ߠ����0�K0��f a���.�%���~V؊��.��,��)���?6y�CF���KǦGixiH�.��S�83�0��dt�v"_���ΙPt��#J5?��$ƨ�zТID������V|�0Z�D�i��@�D��KF���E�ɐ��D�X��_TE��_����C/��d��E���^�R["2����m��Ti�#8i�
�lK���Z���U-����%9�"�@=x�g �t0ě�a
��״TKΉ�a��G��r�;�I@d��^c��{�sp�N?��]Su���1U��=��OXG�P���=�O����G����٪I�R�M�'���\�i�I�����T��7�]��ì06�C����n�: %go��������`d�n*������%�� �f:�mI=��-x�~[�Q��x�{c~B�Fx�'_脇#�N���5��F;_��@�6Y����H�$�!�h.0�\��tL�<���db�j9���{Î������(x��-���
U!G��;�W��T�bg�j���!'T�D@����$�����M����b���I�pj��*�B����$e>eX�;vp7	�(���4z2�K\�x-Z��N���Y��}+�)f�M��?��>P��"�_G��؍}�G���M.�s�Z,�\�-��3��6�xҬq҄��ǵ����vr,a�� ���x5%�r�Pނ��o�*�~L蛒�b�r�-/D����	WGw����I��O�����7'j�p|�eV��Q��Ǐ]�]֗,��Kv#����I^�dU�]�m��-3ڥ�=S��-/e���U�T^w�.^*���/��WM�n�r�;��k�#:ߝ*�vP�B����e�d�[��f/����a���]�mQX���4����V��7����!G��#�]�-ZHh�.;�=����$�HDL�bT_y;�λ�֬�u�ET+�6U�	�
@�:�F���%&a �ȶR&��/���?O��1��Ո�������Th�Ǩ)��4[Y���R_y�Z}�]��?%z��1����Q����3K��lx)��~���sC.�9�I�P�;�m���u���p�@�R�V�4��+G��-��9vq^���3�,���9����U@طRG�g�b��ĴRklg �"Ǭ��<7,SyO#��ݵ���AH�n�%��2�:�A���}���`��h��"�FYQkL��,�uN��t��3i�x@YX�-.�g�z\����fwԎzu���a�Y��=��@�Rh���Q���FF)�^��s��t�D�'�t��M*f7���go���:6$L�^��%ӿO�DC4�}�?9֏U���\�#���`^����	'bcU�ض1�a�s�5�����.�g��D^�@�o���1&�6m�[t:�m�)ޛ�����i{0(�Ǳ1!S;*bdxa̒��ި2���?���V#�^
&��b�����}�a9o��͡�:��[��eL-{�������*ϮI�G`@��E҂��%9�xBŨ���W7�%��>�+k�!�Tc>��]�$8�@�ůƙA�3�~o~Vj�\��o6O
M;)�5Ѿ=�"������I��Y^������w�Fzm*P�4|	o�äW_YÈl'L�d�:���-�[R�������ߢ�-� ��YG9j��>�E&�"G�1AP��1NAHC�ESY�|��f8�sE���}��I�������Um��຺s�C�vv�: �azU�!�c]"�\`��2G�J�:D�t��Du_�d�t��U+�@��D�o�#Yx�������"ǵ��4RW�j�sa+����w���������D�b!����ץ�@`b4�['�W�ۿ�N␖��ȏG}A��Ah���
3�}S���^ �
�WH9E;�:5����+�Q|�Buu:�H�ͼ!3S���(Bp���Պ�O;�X"�g(�D�W����S�
���V������kf�-��u�����qx�����#�L�t� ]�]}���`�������J��7?�����9��^7B}�2a+z7��":�m��.����VH/�F}-E�2ET{}��l=���*�ኍOS.Û���=/���^ҙ����+�g�I�g��{,_��/���ߠ&�G�)�(H/��}�����z )?[��2��c�����N�Z�Ǩ�g��b��◩��[Gy-X��$^���.���E/b�j};N�j�=h� yŬ��z�!g���BX��$_vA��hjq$��0N���&o^>Eo��r�|ٽ�j�'?I�!k��3�%����mRP@���P9v��)��$�;�H���*�����z�0wN
o�z���[F)�\?a���8����=v��@����J#R��JH����M��Ӓmy��-M�!�g�a��r���@�Umc����J�5-�F���跺�����x�EP��T�`Cr�	�Xĵǩ <ͮ�ʫ.�c>�9�	^ B�2��?B˥�~wu��L�[L&�̉7��d=���Smŋ���*L�>+o(`8���ˣ�Og4{���6��X��%�&a��M;�&����L�:ˠ��2v@����] �`Y���%$�� ������Ml�� ���ġ���9�F��<���Y*�E�[�~gPԵ���������u��u˕�@��гP��JI��T���Ԡj��_�:"�w/yK9�����<��M�y-����3���Y��u͕�+~�!�K٬����[:��Z2C^
$DUzzd�a_�� �(Yʐ,A��z��������0'�Ox�V�N� ��~Jp,�&$����G�T�Vp�sy��*/���8��L�����u��v���`�D�=Pa�*�]��,%q��r�@j��+Ŷl�􇠧�ۂ-U$.��
ѷ&��E���w���8c�,�f�x��#�\�eR�.�������UC���ɹ�Iho��^Zc� X�I�8��cɗ(AI7�{r5����d{��	�� 7�6�����7? F$g���ǾW�l�{1F��7�u�C,�V�c�S�D��â�I��"'�2P&dϋ9���}`'oy֛k^�WȜ�JN���J|�$�[@b�dv[�㝆3V�y�x��U�Vg^�eR9�d�u
m�sEV{1��	Q%G�p�7-�{�'S!Y_Vd��{�P$y�+l���d�f��Ҿ���\@��o|���ǜ����p�=�ƾ��bNwM�9�m�N�5�Z�.y�ծ����"��
2��Qn�-���r4�,�0��}�k��OB���Ə��Ԣ_7D	L�	os�5͢��C�\�zb�`U�����K�Š=C���5m<Q�^Z.�S�B_���7�A�1�����6��������М4m��MNc���S�@�;����`dy��E�f�J5O��rkFQ8�7{�]��u�n ���hT�����:��')�2�
/s�Vh�u�w¼�"Pz�C��a�$���l$�B�m��hn��O��EF��҉�JⷩmMA{{2t���.�Z�D����f�6Ffگ��+���h_qw�ܦ#��e�S��Ox���%KYF�H/��%|��d�$���0o�� ճA�P�u+ի?���d=4�A���Q��c���,����\<`ɵ��%qw������}6����U����\a^�I�(UCԼV�|�К �T-45*1}��N�@���p5Z�H���>�����88��~<��~��S�R��	q����-A+�*�����V�E�͟b�at��
������	�.<z��U������m�쓽�<��1x��`Y��U�.���6�ת���� 6��R�UC 8�@癧�ڲ����'��?�
%`V�弬����&��:hi�쑙g�&����;�N؜0�33N���ڧ�Q��WXA�8J!�oH.�\9��K��4D��|��N~#����b�D>5��o�O��(Ɍj�>�N�(��5��o���Z-�N˒�oJ� *���e��� 9�Y�/Nb�����6/�u�cd�?�W�����]��Gì��[
�/�����N��%p	w$t���)�*p� B�f{�����Ȃ�)��Ar�Ǡb{�T��Zh@N#��*���!eo�ַ��3vH�ί7��m����-Q`�#sZ&�f�7�}g`y �&�d!?T>æcΡ�_z$���U�[����=�q*������#�9S�P:%Kݛx,��Ej����iڝ�@���{�B�Q.P`8Fyj�h�~�i;���ol��d�sy*�,�N뤏����e���!��|������y=�^���1�
s���r:��4���>Y����@V�Ł��:�|\�4�3����A+�?���F��Zn7�{8��_c�	_;�ox(=ؼ[r=��]ڧr7Ұ���������ej��p.��v��Kt/j���!�+�+P!:�j�� ���k�u����Ӝ�?�l��JW)�C�-9��]}Oo�Թ+1t%�FKnĹ9 �j:$�d���nR/��$�ݤ�(��6CF��`��#�1��j@�U$�R�w��d�u��#Gl�o1�!p��\��K�q"O�BC�؇�uOZ��sW�EןV$g3��+�	^⎇ډ��Ŵ��CT��.��f}� Hʻ=rrI�2�H���Ak��Z9�-d�H�&
h�[��xR�U�V�Ls���dB,�24 ׭d�
��@=���'׿�䠪��i�?��M��َ�^�$y��\�d���ݮ�Uwd"�gط��m�M�KR0®>���ZΜ�J�
�3�dű�������R�b[��^b�z�f�G�?5� e�Y�n�#-��\]-�Df��*�	�?:X��'~i����gHƗk���u�Ci (O����D�#*F��?Alf���C�lj]��8B�'��)���Ւ,�U��Hy4��	���A?���I�2�w��Xg��M��0/��۳�������|aY'-����TG�#�f��]���9O�Q#�N��JK��m��ʝ��_'#���f�2$��F�b{�DQV��J`�c)�/8N#&������ܨ�aO��;xNr���PL��n�~����}�}=̽�Bj��'|L��{�m��:����%-��@�=��������K����hKf����K,���tZH8�f#žA�a�@�ݚ���m�n�=q2C���| D�My�_ߤ�����e����Sk�+��mj�q78�Q��,��rC����m��ڳH"�I��N�wݥ��@�zm��'c#ڔ5��8�����Ls�s���4d���/�B��aD2�&���.p���&�I���]���#vc���-�~E�u��OA����i�$>{�{:|"��h�p/����6���m]�oG���}���R���V�����5�B�GU��ת����3u
�~��!���Q2)��o/����	
������V�i�_wb˚�J��m�v{��c�&��A%�%Q�Y�B?��m�C!L���+<�^���%;w\;o��*��G֭ۯ/1s؉'+�"��₦��>#��V�p��k�E���ü��
[���hC��o�v����*�XF;˾!��`��d�+�E��Y�ގp+��H{�2��	����c�%������'�]D3��p.��'�L�[f����]���z�:*���w=�J�-���K#%���gW���p�C��{}o?�[�L��>'M"���P6	���%jz5D�\e���k(�����
5RG-��:���[>��d�ư���W0S�����<B��Z�X���J�X-��s羚͡\�P`b�����z}U�0���(����<	T�^}�)������ou6x0j��3������$��SC�5���V�%;=+&�#���Y���@z�"F&���`���<��}��WEʬ�o��|��&����#p�3�LN�*-��,�WdJ�}�ns����i���4���g�����=�2+����)>�|�:��7P��֟�l$�X3������d�e�_f<����`>ȁ<�ba�I?Ƭd���H�~�`�)`W�:ҹ�v{����\�S��p��4��l��8��-��ף�w6x��a��r�f�߿�������n���nP]2����}��슜ӄ�
r�����~�=��<�m��u�؇��.2ׅ�ޢ�k�I��5=������U���LF�/`#d>{�CS�_%�[�H�j.�;Z��W2~6+�[��ʎy^�s�F�{�Ւ��FWI���d�J���ƿ2�G�	L&��5&��Y
�hS��چ[����+���KU#'��I�G�F_Ơ����zj��w�I'f��G�o��d��� ;I�m����U3_���� !\|��wl/��2��FO	b*ߕ�^��\�5�?�P�����K9���Z�1|�S��[Kz?����r˴O.�P��2�%tw(k���c��}�z��%h�0�^�5�i�F��xu�g�I.*�])���Q�0A(���/��h���iڋ��YD��^�^��闲�əR0�eQ��<� {i����!���z\�_�N�RʲkH&�4Q鍁xo��������4�^,ZX<x	��|� �+٠m����+�Pxℱ��0,�l��|�7�����ϧ���pi��6���_�B!��:��(&�b��[�4D~��X� ��ߚ��V+�0����f��*��Z�^�J"l����i�!̆��0�1�B-���슀��']>;d�ă%��\��&;i�h���sac_s���gD;��h��]��;��b�WT�6��·��0>��`o��i��t�5�wM�T��V���砇�*���9Zҭ	����^-���i1��.�D�X4:�.燊Z�2Z��.u��wJ�R�も�d�2fވ�(V��Z̈́w�R�v aU>(������Bƞ��r��}���̍oh��r�HY����Dx�����^��TB<^�a�\��Q�]���.T��r��2:*.oј�?W���?2Ŧ��}fΠW;ঈd'�z�A���,��fQ��!���� ٭e�za{Q��|��7rVl�J�s�q�t*�wB�n&iS68˭��p��A�s�&ڐ�rQ=�y&��,�z:�ޣ>�T�D���^P�!���`��A�A豐�8"%�G�?��w& ��:kV@��
�F� ������(���TG�nuqs�7��Z�����?�E{�����ҡ" U�x�KF3���MQ����h��߆9OX��J&v!�t�k(n��8�fU�������_�+���̽��gV��z�'X4�ZxOw r*
Ə����P!���!�t|-P��~X9�>�2#�n	�wm����hܺ���]�x<n���KW��E��j[�O��s�8"h���w��#i�	�{��5Q�YH&0rm=�}`��+8n�*RO������˽�S���\�6|��u� �g�D����+�P��V�����4�*S��	"��D�%��҇3ɆB��f�A� ���g�|6��!��lg����L�^a�G�1N7�u��&����1���\����h�Ӝ!�d.���0�D����.�=���g��9���>� jٴ���=���v7A����\"��$�5kݢB�p:����ruM�%:����T��8����G���ĕ�k,%�2~gq�_�{��Gv��y������O\u�!?w�p1g��6r��@�=�5������f�*�>����B1V}g`|cuĔCnM�b{�W�m�jފ9��Y-q��cMr������MF��*J�����io=��1=��M��̟��UdS$��K�z)���ZX�t|[b��p��?	[�9�ڃ��
Z!�c���m0�H��O�v$��9"�r��vI\�EzU��p�5��59{]TjxJܪ�Ө�oAS-�3��V_��Y6xv�c?�>.V�{x�ڂ�Zպ����2Q��iF��#��2ѻ|����4�7��$As���]��xMT�\��Uxe�iI�0�|�8v�g�7D�C��&ܠ�v\ל����BZ��J��9*�-O����ї�J��웨��z���QOA6|�q�:m���2��J,�ȰB�{ݩ6:�ڂ� �`�Ѹ#�W0�$6��[p5�'�̉�Y�?R��"z��0�J����G�C����M�	� �|�y{��� �T��|Z�����L|�]p +5�COHˆ�W�����B��Oɴ���pY���[Tn$��Hl�;����V������CBm��6(�GL��h�0��;v�UI�bda��uNC��P�~|�eHHH%�X(��t5Ʉ���ep/��1<8�fؗ�R���.̌H���nߕ�^{�:G�5(ԷS�N�l�+����Ic���L�����:��z�R>��<*`��:�F� �&�,��=$��F��)#v>�#���v�.�熈���xde=��Ǫ2�k��i�����3
�e�l��t@�S�~b ���i���������g����d�g�7��3���xI�4��Ekc!e�d��I��؉r�=���Clj��BS�kud�fp��7�r'1���a$����ł����fq袲�\2q��&5���;�pn�wC�Lp�<V�y�����2j��/��g�:�K��^�YJ��Q��u/�(F��+:�
�
���5|���t��=-�Z�Fx����"r1u!��u�*��U�39sK�D֢՘�2��"Fy������� ~�?+�r'�6\{�t�o�G�KPTk��]��&�)�\�s�8Fn�{0=�J�V�\�ܟ�=D�A��R�b��!�H8(�Q*:.��RT� ����3�m��g�C����q2@m5�A��p ��2�I��l<D���ث��ON��+5'�~�,�������tdDYy�V*��:��1l:��/�r,��� �aA���ݹ_צ��ݴp��b�P3�v���:���uRB��]$�-���	�*2��}��C[Z�G �k���l��t��c����>j�W�Pwp�6s��`�F�4;R�DV0���ra���$�A�`tDMb����m?ȋ���Ʋ֥pU1PV&�[�%P�^��o���?�+]�	�����v'�ƶh؇U�B�h*<��$ $����m��H�ضP��^�}'�.ALZ�����&�}�nj)�VR���p� ��Ms7����r�le�Z�N������<��G?����B�{�ǽ�|Tz�e1ټNO27=�:�6ƅsl���v).�+��h'|c��@��Q�Ʉ��T쯵��s���E�2S��@����i@e-�����m[���2���<���w��f�$���ARoV�/�;��6��޽�'�;��@����^�f�"5�ױ�py��g�����VF�M�40�E/lPkK��"�A|Dп�e�Z���'�d�u'�0�"5�`T�P���B����Fu1(7mdzE�<���� i���[l�}e���k��0���1=�;�DDo�G�Qoy\��ޠ�?P�&[ȇ[�=���<Sxg,,s�ft$OZ�`�}+�-��`�RG��'v�f��gx|�����V뤬A�#�.A�>��L#i�%����k?��Od!ۑ�g�z`Rc=棅��c��]G#�3�Ex�ϫ��$qu���u��T;F���t�b��7Zd0�����-8AbT�P���}�����r �q톚Иy��\���'{�dѦ5���F#������V��	��&@?>�� \�>��_�CfAC�DӮ��Cև ��nBae�����(�M��BZ�0k�89�9�2����R�� �'L�3v������:���;��Ap(�ZT���7m,�1j�i����BX��s5�,q=����m�P;�ͥ2r��+.��ީ��J��c���F��v����@���*����*Ô�� ��v��)��y�q��>@
GR7���1�W���кr#�O�^�[X Lhn5'���쉼���
������������7��a�r^9�oe��i��^5L9�,!���� �Fe܇u�)�,/��菖�t�/��W�Z������׬��?��N:���u�C��+>�5��Cw�9� ��*R��;�[�R��	��1:TngBë,&�a �5h�Ƅ�/��T���&�[Lց`0Ε<�_5�P����j�4d�ND�i�����`���F1/$xN&'�d=A-*�����*��]�i��1��<���0�cy<��K��+�?$��+������Pmrw�Ҵ�09�!!�bu��Z>��X/-�陧�ֆ�����9�aN������c����T�e]4���Me��̊��Dɤ�	jPff�H9��ɕ��ԦUN�ɟ�δA6��y"��T�d�Jł��bxZ݄S��œAޯ5��Z� ^m���.LK:�Z��Kzx����Ǉ��/*�T���f��*��f�j�����c��2�q��)���}�j3���a��?��� k(��Xc�F����2Sz������KR��9ƴ�]�̠�>�hN�7�*?/�q$!��A�v��35���Q;֎}�N!gs��倱^�+\E�[�h��Z�қ���`�s/�����u�������Ls0^J������8�7R���-]�z��:���x�Ö���)�$���F�d��1���a��u�I�Xn��q�0�`?��Q��CI�&ERl��6f�?W?m�s]
�����!���l�?~�Q�7����������7^s/_פ�w�v`{�;>���w�G�S��[�u��"U��>
�W�;��Lv�Wv�8���<�Om&Aۈ"ʹY�*$�B.
	Q&�Tg��Ӑr�pI"�ո��.�(�x�����Z_ED�&�q����l�:�v��M���-F�9ǻ�_��Kj�g ���:����ڜ��Ps�k"�|�b�� $��ے2XNN�dV����6�HhҴ�B!ff�x�05p<�⏢ݯۙ�}���������A`����MZ����	��������U�vK�;�)`F��S2�x}4&0�6�����&Vj&UψĤ�ݒ鹑D��j`v��A��!+lݲG$F٢p!��]��;\��<8i�rw��/cC�֊�|!����il������|�si�fZ��m�Rٓ��^f�C,V��O�V�8:�"�VC�j�h��
�g����g%!�hCBԧ<��V�08ݵKQԲc����������a�����ʾMJ�g7���7�Ҟ$j�����o������G$���U��0ˆs�\�D����P�T�S��[(�9��س�M(n�w%��C��r�:xU�G�j-�c�/���~Ѧ�]6�6kyv�׃4��,����|A�N��8%���:
��;V�M�`����@,Z���՛�BQ��X����-�K�=x$�P�}'��Z�a�����g�=�p��ږ"�w�rj'���� `�)wOI��p����v�嶊e�6|	��R�;�C��z���A�r�0>?lzR���k��KSp=""A]57k)5�6�AT��(o"�$�\�����g��m�@����gH�Ѕ`@�kh2�@�ß ��MU��q`#s�<�y!)����Y�Q[�2(�YN�OP(;�g�\��(nV:�=TcJd)x~�ԅl����˝�mQ����2�vv��Y�����rW��"8�Xq�V~��˞��]`�<k�����)(�ZJ��x�5H�0�gW{��^�=�?y��'�Ů��K�'�L�Y��<Nm@�qE�'o�n�z��a�gM4�����b���Q���u��� �g�����|9 �ix&�3���
ē�������t��8�$�Ө�qsꗜ�)O��^��G���U܊|�{՟�_�d�?�揥l^�4�9�d�#+ ��m���l���ˋ�Ic�B�|�T��$Zk��$�Ӝ+�ߌB|�|c���c��˷<�l%����N*���)(�L�G��� �G�q��Q�EIP���$�^.���8~�>�e��5����ƖN��-�GA�ǣ��	��*~B�ۥJKy:��g'�3e�Z(���oV3��NX<��ѭ[���B��/�$5 ���j�W ���x�Q���S��Ts��ڀe .����̘r�ń�._����J�5	rFY�:w��|O��ү�z�g}�c��Q5ҫ�`���:&��P˻"MQ�!0,"S=b��I��'��rc�r�g�*��n�q��@�$g�g���^^���S���e�>8S��Z�T,�\ܥ�EI)�[ښ�K.�������/�f�<���{���[�7����O�t�}En�7��(�Qï���gfɌ��i�����g��;�����NX��OP>��ōP�)f��/d��;8�N��Ji�q���,Xz��vv�ݣ����7ͳ���XN�n��!I���5�H��yM�ͫr$��n�@)�[��/6��ҝ@��H+�"|��C����2OCc��X��{f�N�`l�Qe�4�W���!i��4�Q�حK���\��|�oF�XE���B��	�B�2W&6�	O��PI[>N�6��^��j��m�d��nA雓1�����Z<���F���C�����nb��m���FKZ����RO�B���2�晄�Y��+��0�W�Q� D|nBT��:|4�[ ��ޅ2!OӜ�ȫh�����.3-�L�R���p=��UP���;����1�v���I�H����uJh[
��Y`�ʨ�Y��'���݀`Ҋ�8T�s���7s;�{��l)<�VN�p��Ǝ�ts�)�_�!��sE^4����I��oJ�+̯�=�^�3S�xޞ�1ƍ��3���T�e��f�s��jO�1��q�C��*�]9����O;�6�y1�\L�t�vbJ���O�]���%%L�	�[|N)|�����>����|2�7U칖�-�b�;�u����s���Hu��)�Km�r-;�|�*Z�x
F��Չa%~k|)pD��9�5Co40 W�_'��g?�M�P��>�x���9�������dm�Sv��N���F���h�޼��@��V�=#- �������Z��;�ȇ@��]쾮� ������BSN���ϔ���z"m��6Ms�. $� �=�xE�1����F��Y��~ ��_�˳;���ɇ�b��ڒ ����4Ūi�`.ZhmV�[����jJ�6�^^n��)$���Ѝ���K�R]�3\&���� ߧs`�뀮L��JL�jrwU"O.�d8�-C�����%s|+e�s'�T��8ރ相�k,����*�{_�Ϥ��-7������=r4.$��z�R�Ӌ�oh��n��S@+:@��ֱt���8���*���+����rv����L�C��Z*�Nߪ��݋�t��;r �]4�T�~a�^ct�)��o=a�a������ի�h�h��ǭ4����X9��?��ˏT��*�!�u
Bؓl�$��IFo � Ϊ�Ρ�hFP���*��a�������5�zu���'
��6����Vt.k��T_�XCܢ���=!-t�jv8A��8�Z�4<-��k�r��w��N`�"˫*қ�<;'�&�[r	��C�A҆kr� �DZ����]�����N}�7pe-s�Fc����L?yP�(�P��D����U���{�#�hO�U�=%J5Җ����lE���x7xM����؁�m_t�ಷ�O����>����n��U��m�׾\�N�H�߷�a}˸A8�>Y+�����T�ɾ��i�|����U�͕ʬd棂G:3��Pln0��M�%V<�
44�*M�e��	}���o�;G�����%0��$�m�/+���p���0r��Q3�P�x7�	l�^4h��l`�֢p�S#.�Q36��#�DU($=%?+��'�ìo7�a����Ѕ�g��)o\ ����A+�����"�i�AK7��n����%��L%K�}��6�L���bDL)�>�����=���߰j?�	h���zdH��Ip�q!�wGŴ�_�\ �n�����X�,x�5fy��^��G>&�v��1Z9iOI,�M91Ǧ���轻h���ʫ�J��{J�	¡�������'ò�B�x��z{`��H�Ϟ�JR��DK�A�1]$��Q0� a��c�Q��'�=��g̱{��8	�l���Pr��������7<���KX�/e*����j�����|֫�5��h�e��+ӓ�v��SfIH��\b=7pu���r0�į���2G�:���V�%�T[�����&Qg���h��[VZ�{� Q_w��P�	���\��M�� �ׄ�L�o��1�3�
���&�v��BO�����g��EG�*O�p�^��S�(xi��B$��&`�M��:��V�a,��/��k����׼(��b4{ᅽ�J�^��x�g��=�3r����4@�[x(�3�=�0pUR�D���\�NGp1��r���q���nms�A�o->5YRc��U�]���7;��7E?aP(�r�a���N�����\|A�G�U��M�w�#�")S��`�U����4[�6��o`dlg�H���lI*%�j�z����9��C�C����� ?�%�!w}����<�P�
��[�� ��-�ޘZ���؊M�3˓<`X���!S��r�:sey��*��j�M���\�w+[��	����15���Ѧ
�5v +i�CYϚ�/� 5$�W�Pt%V99��%Ez2.�"�q�+կTN]���cku��V���습H�m<�M�䘦�PŎ�&��B�|=O7~mc>�ҹ�}�ϝ�J�����=6�W����E��t%�ތ����Ĕ�T�sw�B�cRv8Ko�	��Q};�d���δ��e��J"}7���Y*"�B΂�Uh�o�����:(� �}"7C���m�!��[�fQ��a�x(���W�Z��.��kFd�W'E?h&'��"Q�����̹�v��}�_�-^� ��}�N�C��ptU�`�va����3�X�`�<1^1U)�1X*��v���D`bNnd��,KRX�ꢔt%�z5��]�ſ�V�EWd%��x��z�*Eʚ3�H�ҕ���|u���;�a}�������!gP��mq�yiꊄ��5ō�fm��.��BS��ER�������;�hT�k�-;5�'���������MX%'�`���2�`Y���UG��L�`�M�Z98�o�Hd�s�-���fr�;�Ⓢ�P���w�j�⥠�Y`�b��9�0Dxr��#�_�'/��,�}�`zA��iO���M�[��pj���`�M����:q?��2���>�CeG�bG���V&'R�P�UK�6����p�p��$!�0������FI'��f敘�������t����W�;r|��a���L��V����,���A%�0���B��*�ۗ�V��7Z��
r���MA{�ɣ�W��ʝ�.�s�΢az��_��ȑ�)s����.|eQ��h_�D�A��m��׷����E�jP)��B&�Y��O)�����#���O9#���H$o��Nr��)!n��ɫJ�Sw�h�%�d�;P��!���pMJ��@=�=4��\þ��S2}ܕэ1gL��bMR�{đ;�%��ٸ=��B�c���hS��;��RڔU��5�>���꠮bQ_�.�d���F�wUB\]�8���έ(o�_eG<��Ih���L�.��v��(E5p��D����E�Nç#j�J�P�s�m��n�V;�Q>�V�}���~�#��HfdA�T0aQ����O*���҄y`�Z�J�MZ/-e.`$���-�kN(�\m9�d���i��5�k*v���!c��s���ȫ��$JL�e��]g�	��x6$B�i	^�;LFK��>�O��k����#/�����T��7u?6
��+tŇ��G"_��1/�y��B0V�����ْF�BD6�kye�O/a(р+1��G�xE=����Vj���B�9+$�ۛ�<�$$a�El���g�S°��u]���� N'0��vwb]� x+kj׭S C�0�z}�����m	鯛�s赝X.�MgQ�S��I�~}/���%���~��h��]��X��Ҥ4_��k����R�kz!��;��|G������L3Fϙ-������=�N���W1�g��/����"��=ή!z��
l�&�!�Li��	�X��<�GW�η"��6H���_�P�%��p�[���0@h��n�fx�&d8����<"�^bI	�L�}K��K�-px9���$�r��5.b�����mJ�Y�c�!U��҃f��~_��/x��W)�ŵ��+n>D�o~#���7�а9�5�˕�*�(#=���R[�����.�|j�q����JF�2rVL鄨 �jԠ����)?��Fh���D��k����!�	Ab��|ȅ�'v��B���_F�]Z�
��lL*�`H�,�
��/��i���6���q%��ndE��hImB���u��m�*}&��X���ph���l"U՘?�Q.��Tq��`��2&(c]+f{�1l�#N���O)�.�3�ѧ��"J�����N���J�R}���#7��#Pg�evxH"� ����Ld�"x�j7]�Bq��[(z�I��k��Os�n����ʩ~+qIw�<y'}�L��V�Du+�>�������_�;��]7�������%�W��osZ��9Q�N��:�#�Ԑ���nb����=%��f���(�(�cZ�[���C�,��ktY>�mф`�y^�#�TG�E?}�H�]XB� ��
e���7s��/�2�8�fgҺ�𭸖���J��F!ŉ=�}�/���ҫ���K��0!
�7b�����k���_�-�I���4!y���������8oM��U!!�X�W䭇�a.�h�4$��Z�CX�c�V���:�u�k�}e=E��?��?��X�u��9������������i�:�@�W)�t��'����}#a�]��PO�<���Jǒ'Ae,IR��7��ho����I��pE�vU� �+�P��w��L#`�&��\��=�߻���P�N�~�Ϻ�a���E���]ɞZo�4\��ncls�4�+�7t��;�f
���;ν_���?x�(*}�na
1PT�M�}Pq����c���{G�4pg_,Fä_:�b��2c�����7�U:�h�&�YW�|d%Ӂ����;V����>W�&�.��v���P8g;�9����*�xW�p��d.�N5���Yf[>W�p܎a�$K~��x~�5 ��VOl&�3w��1�;{���0M���N����!p@�~W4
8'P�D�=�����/%^�mD�`�V_�z�ȅ0@�"TI��2��ZD��~�(u�w9��X�y�?�5"�c��R K���͢�%�/f��SZ2�M¹ȥ��;�������6 }�@�òS�+�5��
������RRD�)p��+~��UN�VyF������K۽:���H�!ݬ@��{PBIiZ�pr:�bAi�����o�mD��C�,�f����I�\X	�w�M�F,��(������G_������6p���	�g�d��oW��6;�	E��4�rC7�=4t&I\�p?)����ɛ��o�qI����;�#�����9�|�&��*)U����;�)��	���ԗ�Av�-O4����\Goa�[wt���)_I�q�DHP�q6��Ət�ǉ�v�����.�.087����jt�Rh�̎���X������x����x�3�\���0m.(lF����s����E@8|<��h j��*�kU�(R�0_6�@�A4]w��sW��ݨd!j��]�lǔ~hRP0����0� ���҃��S���x���:{.���{�75�U;2�"�� �Lv���zC�R����� u[��fcX#b>Y��_���M��L�q{�8�e��z�璦��@EcVP��z"�@<Ye����`�ZI�:�z� 8��൞Mפv�
*��#���������N[�b{�dw^��#��S@���Fs>���Wp��>��D,��=#}vy�վX69��75�e���?J16�fh\�����w�.��iF�{��v������0�܉���JA��oes�3rV53ݚz��hR�O��ov&��BbYhh�lj��eV�k�Sg���4��U-��ԒટUNS���Q\��B�� ����	��a�n�Ey���9p~ �H�_��3�fS����s��,s)�+�����d�R�ϧt���$�O����~]iym��gQ�O��o� p�8[Lt��&��%�|�̛4�Y{��Ą0�d�A�85�DP��dQ�R�!�<�A�n�T!�8�B�45p��@�g�QQ��V�&
��a0)=�S�!`����vfgp�(R,5%����I�β\\���Jڐ��*V��1��eBLm������aKJ�b�u�������=~P��VJT��ٚ�uwk�����_4�t?�S�����J�77?9a�_Y8[6��1RJ�|l��8��۝}� d���R,�+~玽�!�c�'̪�/���)^(�f����ì�#�9�V!>�q-_?�h:�@�����Am�`)�8m���c��m��5�V�1y��_����O���T��X���v���wd��N�j�z������wY�t҅�g�A|��K��ɇ���u�����W ��s�?�[�_g�!�V�4�<��c4zO�v7$��$���b���,y����eF8�kk��;�՘H��|�
%g��(YnA
MܴaEk��0���H�+�ƱP���SA���b�~�T	�BD.۠���X<��DCf�?<�;c�+H?m����s�S��#�K<����'"`��|��/5����M�6����.-���+-5/�|���"8: �.?%�x�~c�SɄٚf������\�p�����w+�ZsJ�p �$+��w��|N �L.|����NenLͣ�'R�����!��䭔ϟ�b^o��N���@5���Ba���A����"�"m���1;�D^��@�$�WRx{¡9m�ﰘ�JG:�W���H>����~{���<Ӈ�v��'^?b&�k(�[j\���u?Ňk7%B�l�4+`���T2�v��9~�P���'�ǰ�o�e1�;�����c���7;�dP��D��Jź	P�3\#v���JU@!���i:�]�5
����7�a��3S�1�/�iä�*�4^LA�����k�h�O�DhRM�
�@#΁���kp���l��N�E�H�x��^T�S
�������+�� W��TI��u�zqFU�*,8�Xe���S�բ|���w�'��\ԖikX+�I��ކE+�n�DѨ\��	�7�[�~mr�h�ҹ�M����2֠��jrjX�V��V$f�9��<~c�y@`�c�LGN�Y��L�G�au���n�ィ�7�Z���h�3�;�L0LJ�Y$F4�g���NtJd\���1��V-3k�.	��#q���=s��{����d�����W��-� ����`n��)����7�ۦ���JW ���Ù���t���z�<��l
C�����ᣝ�,EQa��3t�25E�	��E-�r�$�#�SذO��'����:�p���-����z��i�|~�]���&xtW�!8T�u�*P��B�ze�(��T2��X�/�ӽ�{H�JlV���N���S ��*C������0��*xu	ʊ��'>�����a��I��{��>��z�Ւ2�w�M��U�7`~�xF���}ka�4��{�Y�+���M��6�o5T��8�$� ����	��H׏�HCG��72 40��4�$?9�:��$P���"���ƯE2��E���L[e��T�)�_�\�	�Sd픉- �5b�E�Գ������uq$���!��y��܃MJ�/�~�f��'A�ޜ¯`�O �u
�#���g?��,�T����g.�Z��S��O~σ�� ��6?^lc>�� ����ZJƢDt��.�=�|=�$W�7Jy��3ʌ�X�oY��"�=X9v�f���a����N���a���m$����;����4�ӛ̺�?j�MX��5�A�����.��&o�B '��%�� ���Y���K�y��ʪ�^ʖ5_�H�)��
*�?g�?�$W������A����5l�dS�fc�*�P�-ՖdZ�,>k���i��+�ġ�΂�@���֛����r6�H��Qj.�I�L��"�g���̠WUj AeN�a;��pH|ˁH�@;��3��{�W�]|�E2�T{�B�i��i-�����|kb*۪�W�=�ܻ���n}��
<
�0�&�Y�ƚ�((�/T�^��V�e���Zh[{[
��a�s&,	B�Ͳ�FW��ǔ1�)2ɒ`��m���� 	p"��!Q��,�0B�`I�i��0�{�k�4�2JAK*���g�A$W6ʂD$wŶ���G���I�(�ʮ+f�,3Mk�V�k�,*�4�	DHyc�	R;��v]=	ǁ,u��ب���ܪ�K�G	�)uQ�&��<D�U�H����pQ�A
�:,��ς�����%���0�jh��,H2ɼ ���/�o�%��P�yJ��\ǽF��X�M��^IA�QL"j������a���Pi�c��m@bp����m����E���HZ�^��T܏�~�^�����e��/��k�>y���NеrT'冲���[�����\�h���g�cL��Twu:O����T ֕� ��W�r���J-Kqb���c��!�?��j�E [l�1��,��P4��,M��Z��\ʵ	�]ƌW$���yҼ`V����X���*){�_�$�z̔%��y<����{$Dt���Q��?o��܋͈iC�fx��<�Th����.H!���_|´<��'�|4^y�1�F��}۲�hЪ\)�5���o�u�W~�A���9yQ����ۄ�7|:C� .���F�H�s���π�Y��5(�2c%^ඁXEJ��&��¶����Yl�ഗl\I�T��U��g�Ԯ�y������{�R����45�)-�1/�Z��>���N���=���#:�+�d�������5���Z�E�YA�
煪��=��Jab����*(����k�H3HRI�v;/��k\� �̊���`��}ٵN��}�O䛌n��N���Aď������k�x��f�nY_'��2%����*�%2�.0X���cۗL�\hh�n3�Д;G�Iua����=�^L}��)v�f����32(j�G?��\����ͩ�%�?w�G0)lq��uցd��ͦ4�Nl�����Տ0��������pd�i�h�cZ�v+��@��q��Max#"��p�VZ^�9E�Q�-�8�W���Ar����M�q�����9}'E�B8����Si���㐴�ݪ�b�s6�/s/�����8��S��з�/��-�qtU3����y��?l��MJ&ƮZ��@��榋�d�����|ǁ���6�n�?`
ƭ���e���x�2V�b���F�	� 3<���ߖL��^&�b�f,���9�Фl8�����vz�É�~�����f���zd��
v*tc�W@��?O%�����7s��K{Lu��]�<ċ����Y�^:���%�H�g����1�{��[u����S�HI���.���DZ�u����1���*dw����ŉϟ�+�^t%�"g�uA����/A(��ƒݮ�r߽+�*kN➃��ͮ���i�Y"�=�gH���J�|eKk���O�9y.�m��ݾw'=V�"���p�>Ϻ����f�~����5]�ع�,z|y^Y�	P䄑g���AX����A���@Mte�=x���Nɡ�Vp\�p8��Z)��)��G`� ��)&�<�X� y��������ux��/�3�i����zЏ7@�z���͔uO|�)�3q<Ze�t��j�G2Ut���&�� �̴�=+�����I��	 ���{]o����51?]��ŷW\	����Z��Κ4�s���M��P��%@	p���\X�؂\��Q�
���2��HSۡB��٧�f��pJ�p���UX'��V��8}�P7��)⏝rǏ�9]����%@�;u�AsXg^"��mO涱R�-�2�	'e1�/&����1�����kb�i�_�����r8�Bw��n(����eYll�ă����A	}�n~k���y�O��KpN}�T���ɼ��
��.(�����!��N�3hf,Z��+����^;^'�A"��k���3K�Q���W�	inkDS�3_�Ơ�%?�1�wŋ
��庪2:Ҍ�ɟ��7[�R_\59#��Rt}��{�4T~*den���Z�H|�����
�?��Eb�ЀƤ���,�˟8d}̄�x޾�C\z��f��e���ƻ����-��,;�� �PS��)�x ���}wWS��
Ĕ	YUBk�	�եgᆄ��ְ�(�Z`�h�u,��.�d���I��^o ��M%EDAu�W�ˡ���Jņ�As���<?�\~BO��\��3���S�DC�;�K��Q,e	���mw� �_5�|ƣ��Jp�0���X�=�4��z'�nRV��'�p����z���Q-C��9�(��}J!UB���Z�[~q���#PA]�mA��>�''sSo��������x׵��9#t9���+�R6Տ;�el�@�^omd�4H�JM3��F�⡢�t�4�*���0�t��,5Ԙya�p��g��[��cJq��d��d�V�G��{��
�؛��9� �'��O>�{dZ�QHȝ�G�Fr�@�s0Uk�"T�|�{���~����݈�I��r����ne���6B҈S{��5�����w1�3r��Con�\�XL��Lb��%X�	Glwߺ�t�GѲ���2�<����|Bj�H������ \�q|$_�[:)�u����2�է��i%͎� L�̲߽�,�ʱ�Q겞:��(��:������F���.|�W�0f=]� ���7|�H�/n����|J�y�8��s���d}�np^��|`(�)�^簧��[�d�OA\��t紗�O&��C� J ��ah���S�r��5�B9�1O>���������!~R�M1^�����s?6_$p��,�CM/���4+8ԉM(���\��Ց�N������ڶ0옟���������)2!�^{���(�|�"���:'��3b�SH�_	F_��heϼ�hՑz�y��C �g���w��*��cCG�$��,��ˋ��)�('��JM���I�չ � ��7ǒ&���
a1�!R��w>��wp�}NT�dpCR�uy�Gk�������\�b�|��CK�J��x6�,��E@fS����~ڀ-��/�燚���T}�
�����[��á&�|�)��bJ�p3?���r\5�`A��g*�[!5�	Z<\c�餮���O*I'ŉ�KD^�4��{v��όNW`�*v�dbd6���k�2��^�O����:��T�&?=�ػ`�b�'��p�6]f6�=�#�I�|4Eu�bv���o&�=�lb\�:�+:�J���՗��JYh�_�6���|jvC�
����p���n��	<O��0���,�}��$��h�܂�?o����xߊ�������[������f��#�	F�`������h�f31������p���w�`����b{�Q��yyK�Ѱ���@V!���N��I��?�W��v��'{B[�V)ۢ����	��̜ o�򘶿?�RS�[��+?v�R�����7��'�A�#G���B�8Y����q����H����ͽ�u����vd1���	�	�'�얧��!��ȭ�If��� ��a<�E�pFlC�'�T%gƨ���<J`>� ����ߖ�6;�����5u��~!�Z�}�3��(��;l�5�H��Le��yI���奜���0Z�K&�ч�dP5TU�rlkH�Kb���Y��R�*p[�!��!!��Ug�W��pC�e��SD�U�ȃt�5h(�~/4�,����a���y	Ӳ�Gw]S�+'���M���'uh�B�Lf@o{�ɫ��q�nn�����dRL�����}B�_��^"��Q�;|�S���m�a����v$%��o�W���4�x _���3apsT��)~H�Q3w���L�W���f�j�Gt�)ՙ��k�6�?.73�B ����Uz@�^�$ͮ<�Ԗ�Ņ#C�����vҖA��c�[���ح���2e��_*<��[�<}{^=tG9<V֯|��&9��tV�����Y��J���5��W���T_�s�jm��y���[��0�V�<2��'���t�(�=gU��8���)���,5����,Hh���پ�2(���ObK���p:J����J����~��?�'۲ s���� >�9���b�كz�b?����ɒ�Ga9�J�q&D�p���4"�2m|�j��6[���שw�Y�0sR�r�	�d��~"h�����7��(*���zt�<�%���1��٣>W�0���n�B~���=�b�l�!s@����gWsp�[�`�]��X�t]Z�V����`����Ӳ��W����b�V��r?�%�����SY���Mz_y����!���H��孶m�p����c�<�f5{*F�u��������^���jS�(��:�Oֱ\�~�`�d2Б`)Bd��T#���ӷ�	Et>�j:�W ���$ֽ��l�H���QԜ%�����l�3�rU�mD��.�;y@0�U�uo��� �>;����W��)�s;���s:T�m(!Ws�n�,��ڵYWv�C�� ��������'c��U"�f�������e8ԏ.��I������ǶX��O��G�6�R d]�1P��?_��_k7Տ�����m�����`�F�����v���}^\q�F�M�*���	z%�ʌ��Gi6�-�HQg������M�a�K�.80���Q��{J�}�Έ�M5x�G�/�|�mִ����A�$���v�$�Y��t�%[{�{-5��4ba�[�?R��_˗��hj8}iz� �y׆�7ɹݽ{���ˑٕ{ڀS�jfb�����S �5$k�ZE������0(�{"P�+to�Ur==�Y��3���P��2X�u������;Qlnd܄��g������R?F�P�ݷ+婗�`9�YfK Zrᤍ���9Q��*��jGO/fT��C�9J�E�ّ�U�[��G�b�b�p�TF߳[��{�k��\IʻGu�T=L��f3���+�f��S]X&\[��/xo:�{!{/�_:U�F��k�UVqt���!8�)�߸U���X�(�� ohʞ�@��yo�����b�[����#�QJ��.fu$�Lc�y�����v��(&�$W2F�#�]E�7Ty�$�b/^RH�@�v�7cˢ@dS1�$c|�wl�U������P�Ȏ)�)x�g� |�U�+���I��-~�7���Oz��,���0�Je	����h��Uȑ�!�N1��S�`'KP=�U=�a����v!J%%ɶ��`S�^t�c �3���(u��C����lB�(C0;�6s�g����.%�NqG�$�E��>!O|�v���h�.ޔQ�^�
A^�]vF�ĪP����6���������Y(������#�ժ{�)t�=�Z�OydQ��w���7��L$	��-��m(
��hp�i�1\����MQP���Ϥ�q8Z�����a��B�.�3���9a~�dC��]���V߆ws�r �~���2�#��ѱ�$��U�;��/�_x�(��9&;M &����a�/;��c9h#)�zUJ��tg+��O����&�c�3���'��?4�сRv �UX���ۏ7�R�����uК4�m�����i�^�F���V�&5�O5�ڽUқiV��3������p�|��SCK�[k�dS)� Z�yXTBq�Մ�bfb��\^@XͶ�AZ�w����y�nc���7e��5�yU�o��U�p��>uhhc����^z��NV�=����Գ29�����)��Ǟ�͗������݊�����"���\knN��:c�?�-�P�@:�z7y�^��b嫁F���=����4T^i���P5��g�*^�pզ�є����J��k���@i>�c+Q;�}���dCt�7�t�׍Yz�#��r��2��m�3�W=L��=�,�ߴ^�[����+/s5	)jb�u�ߢ���M���0��w��j��NK��q�A�W�m��F��^��({�y�FR}%����^����'P�d�v̛͍5�f�;D�NgL>[�+�2y`�8�����ص&�ܟ�����"�
*i@$Xn"��Е��.s'y���o�ۛ�g�Ih���
0�8��Yٟ�1܍c=��'�o�K��{���gc+�6���@aah�#;,r����
*�;�����⻮�j�'�PV�����I��=!ξFG�"�(��E�䆳2�w~���i�R.��7��Բ."V���u�ʈ�s�����<$��O���7��^���v��r��GD��㿟�h�9����E-���
c؃"E��J�G���Z�������cF�fE�����b��y�^e�ÍeK�HԄ"��i��> ���4g�B+|"Jc�&i�%�0�`��_�IFN[�x�
��u�|h�(q�s&��+�o')l�wϯ0�� 4cD��L�4����J�ځ��R�0�J�޷vl��}� ����E)��5�SýʦCd�\�"3��}ɚr�Q����e@�KZ�{�w���~#HIރ�t kp���u�@�q��䴏fJ����O�_�y���S�"��å7M��7�$��zI�g?}�Ny�Y��K�aO~U��%�� ���F�m��
M쀨j�!0��VOm�����۬OjZY�Xz7�����vL���q��G:�<RMX�J\��˶��t4����ӹ�E�ۢ�Ǚ�d��T��&vm���xN���^�%Q�XDׂ���$�#z�������5k����8l|yji_,�H>_�d,�?�a0�ӷ�t�5�r��ȣ����Q �o�o���/���ƆY�w�%z�"����h�܄]L�0Z&�����C�D5=�H`( �q��q�j��c���uOPQ�m�9����N������5��9~}&���i�B]A��cD�L�*,. �����T��Q�Fp�X���ka"$ww��f��qvn(�1�N��u���7��������f7}���[��g��~mY��)u�C�*��x�T��CW��F��0�٢~e2D�1�^���\򌣰��������?��H�Pno��tڶ��}��]x�o����D-� ����a��G��� l��B�,\��L&��,�軝������E��_�gE?�`��n�hT����]�'n��$�}��=MH�|\g[�y����KJy�Wz���6��Uw�T�W'%��?Y�[�.�j1!�_\K.)*e�K%g��j�_�鹓�	���n���,"_j�����(@g����<q��C��L��}Gi%�0��5 ������	����RZbJ���-g�&���*PT6!yD�K��/a�'��ʼ*1_�L1������ܓ	�.�p�&|�a��醡p�ڴ1ی\b�W�R[E�Uc�Pa������t�	��%ʋ��{�=u#f;��&�$N�>vRs)}2H^���̜�7�G���.V����m���#�
u���'���@N{���3o��D	��vT<=�k�ub�w'���+|	�D%�Xs�W�mi�T�.ψ&dH
��ȼ��"�mn��]�ɱ��7V��JNۛ�s7��n�C����Q�X���E��ݮ���9�G�0�(�'���l?������t9���1�X����sܒ�$���wT��@G1�1����J�p8D������ք�.����5Vo���՘!{��Jx�^[�P�f������ދ�n�_�J����M�C��ʴ�E^R?�3�L(i5,��¤�h(���E���oR�yj ��q�K�f��*�:��3�!ͷ����I�l������Ibm�����a1����E:d-����n�?IQ�Q�w&���s�I/c��G�A��	o����k~U�����"��"��]��b��^{�;�஄rϳ�Ի�>� �V�q��s��Z'͚�z�sV�9�h���*�����.g�2�5�.\Ot��-1?��L%��藩�F���l�ʮ��8o�,V�u�����%�	zC������������Y�B�;Ã��3b�MY�O���%��f��K�����o�a��&.t����}
*G×JC���f�:�ov�MF�~VT��'�]���تA��*Q�b�"�&�X����[u2��9X:��vN/�a��[���\�\"`�G����%���D$E����qߏ�Fe�}[��z��j����X���'����)�k���ݞ�O�·���!$�8��L,�Tm�}6�n+�섫�BS�G�J��s�$�ڿ,���aΝND@��� ���;3C�7�nJ����&�$ג���ԹC	���l�ѫ)^|���"���;{�7'/(�M	o��`�U,���z@�kܜi�x[9��?X���\{�P����ǘ� �~�w*��"6pw���m$E6�n����am}��yœz~� �����1��R�&�|F��0��@��q{ر�V���������\�t]�8�����A,B������d�6�#�@Ȉ��9��p�$Ug.)�B(��"�����8"�0P[v�Uѐa]z�8쮣;���"�-z����@�yV��Xk��5���:�2�d%�	ЃV�õ�g�&��g&�}?r`���0/
\� Ǖ�)�F�X�����V�y9���Ύ6R��X/���ײ���9,y���LT*������Y�d7b�/c`��P����̮�pF�ˆ�|_\�1���U�rX >:]B�q.(|U�底>�:�3�ar�f�'\�=[|@R�wE��V����&�5�D��d$I�G�J����JE�B���c�q�%�#p6/h�;�f�tф����$\ٔ!#`��|W�0Fqb7�� S����S�r�*��5�B�Xl�ɂ�GX+�27Z�#q�%�A���H�\��yG�D#w�M�Y.�-l��n�!�x^� ��'Xe,p�ɘq��>�#�ۑ�Ԫo�f"��>5"�u�,9N&���f�y��U��~�VxƔn��]:"���D�O�[c��+Ɗ�仐E��إߟ$o���۫�� j��	:44`c��~�$g��bIU�x�������w� ��&�����0�&���X~M�\<J����)�!1b��({&�&�U�����⋓�*2��k"D�C�zɟ#R5��L�)������]=]
���o��wK���*l���;�����Ӷ���q~�Go9hɂ1Vҹ������DrX��U9�U�����;�xK'��BD�{r9Y��2 ���;#d�;�����-*x9�O�Z�<ғ���I5���0� ��k��APKjEyp(Y<�\���[Yυ��4�E\<PqL>��A�f��n@M�r�p�eQ A~f|0�������E��(�8����1����<�wҷ{��ݬ7���>o楌��m�M��^L?G��X z2�6 ��F;A���,�lǳ�l��V�x��	�RfC����.uG͇G��O�'���[HN0/��	��z���x`��i�%�� ܆I���ȉ?�g�[�J�S͕�������Dx�'�ϳ5�M�X1��C�o����bmb��E�PF�X�����I4p��V1�����=��V8�+IaEx��*8G����>������28��Y���2t�� //e)5l��5#\�ޠ�-�)��Qy��������`������]��u���U>-���[Pc��K�:�kL�F�Q����{��}�=\L�[J�)
��H)���Dg[���y�F7�&��$��X�����@��A�e[����U��]G�#3�2~�(�%]Z�|QM܌:'{gK�bs������� 0��"�3�`���I��@㉾I�]�b���4Ձ���rZ;�ъ���! q�tT��f��Z�=�y�Q磐p�\�@V^�I�[��A�(�]TpaA<o����M�[���ך7+9���:Lh,g�E:�~�Z����A���՛ݚ!���&2H�b����)�v�������T��r�7���ԙT�Y�.qFj_���� o��yR�\��+Q;�{�kl)R��fD�:G�6^W��o��?��"(��'2�,0�Q�ێ,����m���<Hl�
���Ű	͊�������g�at�"��:��NN&�H�$�g�\�A�9SP˞�O �Ϻ����F���]�d�#�n�!sOU�v}��b�F���T���Օ8�Rp�(Y�ӡ?��A��M�֛Z�h��ʩc��OZ)����		�'�V���97���{@%�Z~\'%���dX;JI�;����DPw{�t;e-���]��ɝn�����A�sح� 9h@�B��wd���t(�H���%�H�/�l;�l�mŒ����O��a~�>�����$���PC�j7�����buP�C�{FE䍊�k�9]O��ZV���%�.ǟ#(:c����o/^�-'+ a �
�.M��F���8N�3����$��<�4G�}��,�pb����7P�������
�i��M#���1/I=g�gb<������kX������,�@���AR���%��9�1�ry�K�R�n�ce���3��U��'�#J�۲q�Uif����%M�k���"2��>1�@[�"b	��Ƽ��+~-<0��Zi�`�\gy�� �L����,�d~K�$ѰRFD��@����b_��v&�y_������D��F���Jƚ�;�t]�^ڡ_s��l8D�7b���Z9"�s3�;<�����Œ���
�kK�F��f$��߯|��#�t�V-�aG�t�����n�����5+gG���dI�q��Lu�P<>'������X��,����{feS q���#u@ֵ�a�PiD��M�X�3ϻ��U�Lp�u":n�|��E.���O*�rd�J��?
Jz�Z=[�/��wG��k��6|xWb�}�礐/a���*���C�������	�������R� `�ts�Œ�W-�f1h	R\ľ��R��+W�c��~��$2�x����P����4�>x���y	VUhk�4<f�A�B�p��D8����$�㙇=�EL/����~���~j\��t[���_E?0z�U	��}��2�cR�w�7��`��f�
���밍u�M�b3LS6N���A<JZQc�=�[Џ{�DUϫz����^�&F��{�ӕiX��	��	��	Ǚ��B�WB����5"��w�<k6H!�Z�x��ҧ�5hܐ�\V��~H3u��0�y���� �9"�|�ѭ�� i`_f~l�؂��Z�5��p��ZICk���p�H�D�a!�U��D�1.GSc��k�`�ē��lX�Y�%^,���5s4.i��:?�;�0a�ɖ8�s���f�r��G�����f�-ُ��aLU�����C������$�I3J�����j�Ϻ�c��lg���#�r �w���)2Sע��$���:��yڷ��U0B����[P�¥��{���z9���
_�Fa~���n&�B��R���5��w�c���4^c\����E��c�~�X4!�%��%Er{�I1���_T��48�2��3L��gȆ�Q�Yf�j�-�L�]���yn�bY�J��1@8Q/���׵%4Ʀ��<�!\f�ya�3��4��g4��{����VY�8no�;�KK{N[�T���¹q�afMbR�ڡ%^]O ��aJ�Y�_G6?Qo����xy<�eB~��yo�9̍���0o$`hj?|;9 C��ű�E��{|���#��A~%D6���B�{܎�c�W#�>���/��9���XU�?Av7�'U���D��J����n��x~�hc�������`yR��xh����pog��i���q�EJYEhJ���#�h#�`�3,�ŉ���C�ԅ���M���N��0Fq�PS]�Vo}���Z=ì<��<�	T��m�ƟO�~2���^��~���#����#���f��,P�U��ٽ G���"�>'-RO�&R�B�r1}�d��� ����L�|:.Rӆ�� Y*�9�d���(I�TӐ�nP��c[����.KW_8J�s$Ӽ0�`1,-��.|�k�����P����/@'Bя�tHx�{����2������/������
R��[^fh"��8o_��1 �z����'�#��J�g������5r��%�8�3�-Mo��JZ�����<c����:�T��5y�$"���U ���N�������qa'���7*	ƽ��tA��
�jKW�����lL�'"��h�Ĉ�'�%8�M;nIv_�i7-�w�`zV����a�|���]�\[ 5�`6x v�#����XlÛ���f/ʴ�ө�D����o�o,���ڵ�������k �	���F�/aU�{/G�b����6�?ۢ�bb��dB!�j��*�)~O&V�}����-=Os�f� C�Y;74��=�T�w* A��M(�hھZv�2�j6z�9�^F����y��SNҨ��U��J��W�XQ�!h��|�KG"Mс�vL�;ӈΉᶷ"��mK��!䝲�X� X�Q\��)�ҵG�
�û�)JWM�4L����֚Z�X�������6��^��[�`���������($!��ڄ��J*��y>6R��m�{H�:���z�U���f��/;��&LTg������Iu���k��L�4�`u
�hB��)(�ނ�[z��چ�)me���t,����aࣔhٌjd9m�^:o������@��[�����Y�a��*��C�J�mL�R�������vz��?�t��gR�҄O��@��Yd(�?g@�W�JFtdn�����+�q&K{���$xc�baAP�&�Yͅ�lFݯdy1!��J9�{\��f��4am2��job��ӌ:��l�x~�����D�(O�%('�"��ӤoZ�W5�ѵ<�=� <܀X*��*�|���V'{�ҡ�N�i�Jd���[D�j��'�h	:t�:�߿V��)���נl�W�6|�O�\{��07���TV~HZ�~��Y��Jޠ�&�nV��iFjv�G�_^ƻ��#��TcB���N�J�ק3n�[ӄվ��FGo�7�ce���`��6���'X�v����n|0g5y�A�%�SZ����$(2]��n
����@�X1$�Z�C���c<�!=-i�J|��B��\�R �g��P�N縜WЛ/�'w�j8w�����W��.ܜQ�_������m]d8��K�U�I��a9�X��[	0�qX�������:��Y�� �[������ζ��B���q4a����9��b�Eh��i.<���d7TC	���6<q�c�r$���A�]^�ڄ,⭉O}©������Ma~�@蝣	�｟HM��}7푢f�`���QR'u��!� �0�WimRfָ�t��T�{K"6�,Ւt���D�u��g�#~:��?�i���8��Ͷ�K��Q��H���&�"����6���<y���v��6���Mc��{]���?���4fR���d�9�r{��M�I TW������ɐj�?��6^�JFۗ�j�:��p���%�3�$�W||ro���Qޝ��o�a��Y��u�Hbk޶�ڒiU�rGU`�K���/	�)⼑h�穳x���5+g��B�����LA�~*j8J�L��(&&\/HT���vi�V�{���[Rc8��lӟ
+(�q��R�E`��i�N(�L�	�<�o-��%
l���Wx;p"���(\2`AT��Ϥ"M��;|�&Ͷ
��ekMu�"������aS+g���VE ������uV��'F��ҍm��?�&�m����L�A�QT%=Ɂ�&�_��(zJ�tz��U�c1Ax�Q(D�2����k�[�j+�X���\h�hT�J��q�}p��hR���l`w:�o<i9��]����\���7U*#������nZ������:�B��:�#n*J�� r�A��{qН'�jb0�WK)��O�'U�m���nzX�����=����к��K+|�`<��If�FAk�D��D�=n}1Hn1��{xfou���`�/��~�%jğ�-%?�t����/���Jhtˤ������y�Qٹ�#s�L.��X�v씝Bzz�RJ#�*`Z����|�:��������������
A?�*DcXvw.�~I]{��;��\���e�����X���H�#>��o�ic��I�G�z���!J��f$�w�
x���6�l@��?L�,���nՒ�:	�
��'�2`F�%t�V
���7�d�i�s[�j�&O�m\
(+{�� r�+r��D�n	;��mMT��9���I�������>�[h7�a��=f*GG���1Z�57WMv{&���T��wXa:������}5]{�9^���8�!���r���Ofd�)k�#5u�Yrn<K_�0�4�{u|{o<�!��A�qE���w\�'� 1�V�׮S�2��~�h�Yx���;]�Ρ�k��Gz ���T��������b���zȴ���cY���	ʥ?�2�)�e)�m��">�����z�g��Ee��q�$�4�!7�%Zr@v`K�nGp)U\~���o^�X+����f�h�i����_X�j`2-,t�I�!o?*4�i�� �܎#~�_Z '�0����E},�6 ^K�8#��]�d�����Z��b9�[�����H�a�F9�*&�A7^O��.�	6�"�^����\d��X�O?=�g��g������Y��t2?���J�W2��3�x��"<�'tve(sG��ih	��GE�G���p��K�:��^0������>JL };`�3�^�<"����+��Õ%\�'������p�H����9��l^���*�����0��	J���cM|�v�#1�w5�1������-׃>�s���O�gjc���ܣv��/� �T�o\<���Mv''��6ҁ�~͜:m�lM�WAf�]�P�%DWk�M�[9��X� �tUp���C�Z�W��L��fٷ�m����(����(`V>@鎞LZ'A����Y	��eP?��"k�T�rtB�'폹.�­�ĠM�T��(���I��	$2��3�Y�!e�U��xr�d5D	�:m3� ���,�F���y��5�qܷ��c�=1����͸2J,N��}w>��ђ�QG�Y4_gWJCB�;�`��$몯����	�'U2�U����ۯ����S��T��1s��{5ݐ<�G�b�/G����o����pn�mV�o-�����
��]҂���/�h���S����uE����;^�{s�ٵ���~J��C���u�h�@�9�,5�8"P�v-��dWVEN��f�c� �w3%(\��+t�A����5��d��w+�g�Y�$� z��8��!����в�v1�=�`ژD�c��mvCQ�tC6����@롶�k�d�����|a�T�A��/�Ā'�2�$�s剾#�[�����(�j�q	"������Ĺ/DdrV �U������d:�,����]��Ǉ��xCt����AAQO�1��b:�<cq�Ջ��or�cP qA�qC�r�������<�D�SGC����'p��v�ĕn����mƹ�35��3H@�gg�i�����ZC��ڞ:�h#��%F�J����E]�N��C�5��kX(�1E0Q�v̕:�O�����$�m4	��%��T@�ft��|~�zlHqh.';�8@+�����D�2�S �'�$kb[A���"����닒�<qk��L��S���  z�eK���z���!l�{�4Q�|����NE�.����wU������lu�rh&�i���Ϛ輚���n��?��P\�a��}��맰�����	S�ʬ�w�LP�.���B�ߝ'�uy���-˰�F���+\L��m�v,�p�5!�ySE^���xa�x�ԑE�R#j�2�U\�/ƫ���D�fl7����NA�v��Ay㺐�M&�y��̯�^@�?�iԸ�b�&(�ԁ�pm9�?������� k�}�Ԣ�mt�ow)֣W�X�ڷ�N�畚�:0��C~�k��I�7��ʟ���:��<b=��`�Mͬ�OD�����{z0_{t7����|(N!�[b{�!��OV�� ԌN~��j��L5�v>����I��m8�H81v�N�� ��
*�0��dr�L���E��dJ&�i@��ϋ��x�gG���_��:��~������*n�IG����zkt̎L�N5x��b�yTk�I=����>O���Q��}��Z)�*��°�+^!'2⤃w������d|+����R�!mrD�Q΢�8�9�,��z�&����(���g���-�SA�o��ع����@I~L̤�{��>�J� ñ
����D%�v}Y?$[�˰�{C���1Wd_[݊s�S6:6��O�X7��6��0(��_RŚi�;���Z�-���2����3х,|�k�X>��2�F����e�/G&Ws4 w�$C��Cj�إ�Zi~���0��D�V�<�a�Ȝ��exݬ"�����+��D����Ҏ>����oJs�B�^���|�7�=��ۡ:��4�Y�v���@h��%d��(	�i1��-`��iD���U��k{�)��b#�ψ�5έ�w���V���Q���<�J��J<�����Xd�
�y���&���8K�=)P��P�u���/[)��i����A��j����y�w��>��F�,���~��m��2���u�\���	�9���_1�&S���ڞ�/'�8�I��G<4�n��i��m�Ml��U:6�����y�"Hh�q�P�/��=�K,��*,�a�oI�k@в�@�|��������i���D����',WO����!>�x5��!J4���5SY5��c������)��5�W���3J�0�IwZU@�/AzAxδ�������n���1[i�Pk��.��+*��m�rt�$�(�׹���o#?_
]i��<p���ѧ�p�U��x\��4�/\��_嶊r+=��4\LI�78�_F���B=��i�B��Wj�X�9K6r1���&�A�w� �n�})�M'�<V�]��+XBu�t���X�0?t杮o^=�2�by�&5	�ȁ�[*GK�\4��^	����7��
���g����.��Wb�9�7>�zwR����UE�c|��$�yÇ�>5�N�\bf��q��(�k��3���󅽲��F9r{�:�#[ .̒��)����Ґ�� 8P"�@��
�|K����
�����J�j���C�UY[�$k���,��r�]� )����UDz|�83����1+�;���8_�z��D8�	����I�d�W#*��%���@���ߚk>=%6!�igxƈ3O�sI\W"��<9�f�AG-���Vçc�'��1�~�#ֶ��[�ow|���SC����4Sk�Y��mA#}p�RC���]�]����$h���j��>���`�4Ǌck�]��_�O1�v~���3?]L5�?Klڋ���h:H~�������[��B]뽏�t�^���*K����}�?/3pɦ*�2Qv�˸�4N��)+�}�yL��[����~��pjZ|ʰ��:���)�6Z�7c�8��F�/�Z���t�}4��X9o�;�lȲ�c�v�hb�5@-�캒V{-z�~<�r��ԁ�⪤�̑x
F�ь3�}B���ʶz�~j5�A&��t ��ރ	�Ǩ�WԐs�Z=n�z�5r� ���덮��$2�H�����7.�)��F���,�f���.�%�=��[����ڗ&i�y�E[��P���s��;�,�S 5 ��PO���6�&�EZd��nV3y���Wl�=��K�[�}|eM�z�w�u���	Z�C�d;A<�;�ȇM������;���������>?ˉ�@���JdӀ|�"Y�s�؞]�~���XO�_��7��?�iF��K6���[$��|��~:橕'Ĉ����F�	D~X����k�X;�4?π�{T����|y~�so�|㵐:��VP��os0k9DUZ�߼�yxoQ�]1(["˞33���M��$�n0'�[��t�N��NE�d7�M��6�g!���9�z�x�;��Ir8�^�d p$`o�]~��Aẋ�~��FY"���3:�n��4 ��L�y'<��9c"�2|��9x.��Km��ғ�A̯��آ�-c�	kM�v�"�-��@@f�CB�Pi�+��l����} ,����u��8����AV2ߨר�ƍ���,�+��B w@ x
rN����لk�B*觛t���� ��z_G��}���?�.L=|��%�M�0L�:��/�����m���E�����PPeXxh�<z��#T�=<f7�Ho��u��?�v����ACq �~~w�����7���"[4Ȥu	cp���yf�������=6������6���߷�C��g.%�_�a@~ U��cBw��H�[Yf��tc	�-��m�.�y���`��V���b���n=�Rl����k��o�cl�z��,e���K�J)$@�3_��	0ONN���#�`Ps5ւ�>���>��;\�8�ͺ;�'β�(�X�M�uklq��	�4(�Etj.03FZ8P�gp�z#א�W�1�D������(�֋�'�a�&|O�G���k�
�jr�ܞ��D~'��Zf(�ҵ�\"LB�������Y//�@�*%q|�˗|8q/�_Q�dޓJ��:�KVW�1�m]!h����N��-��i��+� <L��-~���d���$�ܤ�-�S9�=��=ȼ�\
�J�5��&�H�7��_]䓝p)�� T�z`�۹,U���i�CJ������W�&vEπ�a���e[�s�-Oq_����?�����
-N�:G�> I�j�lȨ~���*p.Qg�@˯��%Z��;<՘���j�z��<���?I:j\ژ�xUD��;̞`_G�ۜ��R�*��Y]��
y;�1��s��~�u+����Э��<D�NkNԤO��퇃<�Z���~�Cg���p�r&��ӏe�=� �]�ꠀ��(l��8�<�`Hh��d��MV=�.s��v\��ϭ�<�\^��!�(�����RuH�7�v��>�7~Tk��S��:��x����:��Q�vCӺc�#�l٢%�_�R+"��H�X�Z�KB6����i�l2�ןD��/o����T��2�5�0RMB�:S�O����]��V�>Y��~��0u8Dp������1u�oQC2��ZO-�w����9���%v�O�� ��6w��ڨf���C�x=����'�~<�)�yW��9���qe��SfUq�����G�3�b���Z�U�轨�_���}�˗ ����r��d�#V^xJ� �7o�=(���Ö�����v�K��]Id/b�>V��7�	����ߐ��o�p9�Z�O��ʳ��+ kdp�Pu�Z�.��4OK^I���ΞC�O��g����D���%�X7�8IHZ���a㙬��3�A��]��%d�uD΁�Q���D,���*1f�,�ı=��wGpҦ`����V�Yܶ�rܒ��������ݡә�O��+��:�o�kvH�e?P�$��͞?$S�+��n 1�^)q��@aX�Xp��O�	?mU�b��wAjs��2I��T��Æ5F�xԐ$Oo)�f�S��u��>��Pq�G���c���1!tga��ˉ݄�P}8s�x��ocTs�R��~[}���3N&W�#�t!����P�|H��t�]B��V��+H����n(WZX�P:�G��Ų�y��)�8|e2�K0g[�&Ϣl1�5�����
\Z_�3x蜳:�f�8TL��u(뽗(�fH,�9+gR�����j/�X�vr�y�r����o�w
~͢Hv�g�n�<ZN�oLh����8�e4ݾe�������[�8��"�7*�#y��ǟ�L�6I��<�Z�C��K����ŚG�!]*�I�fu��j����	�BG�e}��wn�P5����Y���!���	%x���̊9�ـ�|P��֋ݽ�)"���S]J\s��.�����'��H��	3��#��c#e�Ae�[�V�Хi]IBL��P~��<E�3�~�P�?}�q��
�y�hvN�^�
ק�(�:���V���	��������I��n���2�i {1�@�gx�Z�Mx�7~v�����O�j����X�mŌv�Ĕ�b�f�-�oʨ��/A^���z�k�w��N�rs)I4R"�j�h8�����6<�ڻ���tW��]�k��_����"U#\��cbk%�1�o3#���+q��o�.l7D���7���E���N{SR�[B?+)���;p��k�zG����o��wx_����0ҮC~��҄P��{`�~������ڃ$-q����Ğ�8֔q~o��c�gT�~7��x���B�]@�D=�C�'����E.�V�B�
 �O6�1��X����*j�m[��B�>kq5��/���g�/��k��I��. v��$�n�+��1�J�8=Ry�ǣ~R��Z�j���PW���X�]n8cM&,�3\b��V?p�I6�6c�vll�[Q�<� ����n�:���Ȋs�n�U�Sj�K�+XW|�;"X�5���-�zZ����Y���%�>�S��G7u�m6��x8�r�tv܌(��N�t�N�i_D�9�8��ջ�2���9�W�ˀ��Q��J�5�2���e�L*6t_[�ƾ
W[�pI�����vJ<G��Ix7��:����i:�-�0�*�ug]U�;��*q�� w�<k����`.�(d�f/`bФR.��K���z����*֍\ٽi�x�	�^ky.{A{ݥ�u؄�#'�C�Dɋ�xGD��L����F�Еq��C�9�x���ӛ�娊*��p��]�������,�������T�~.��3�~�.��n��lf縞�I֡�r���2G�����1�r"��J��ԋ�5��Z�ȍ��^4��|��2VU
 (	�E�I�BR��?R�� �a�TDn�vE�sC�
�b�z��.W��ψ�'{�s���v�Y$H����Uޟ:�B��&���܊�4�w�|��4����y�,\��~&�IY%�V9ǖ�cb�^'�#
�@�q};̃C�()��-a޽+n�s�c_�oƪ��j�Z�83?� [����a~���S�f�G�㠜ҭ�٠D��5|��c;$����P�EsuY������̆YT����46��FzE�parC�f��,>�c��]D�6$�f��A�2YoV�OR��<�ϫ�V76��o�Շ�,X���K��e�䯶�ѽ������'�А�w��O��ҩ��yn��B�a���F�~�g��u�o�b��@��~]m��`��c\�Y�H=�� ��&�$J+�;��L�$�n�`�4S�<5��b�)&���`�L#h�v�O����@�sT1UUv���;ɳy�ݍ�{k�z�O?s��ʰE]}�[�%��3�ˬ����]��&P�$������&���Yg{�w`2Y	����Я�'�|Ð�Z(j}���Oi?�-�O�˻s݌C~Y���9T:X뵙� �wH}I���Zw�XU`�\�!󶔈����M%əg�����S�P,�ȗ��m��=�Vܴ� i��߁����*��d�yC��fBC6n�s�Y�!H���[<1�qQ�UoY6��%������3��x��{!���怍z<qX���̑d��F�~�WB#NQ6���m˂q@]�"�ǳlu�Œ�$�_�U�R|�
�P�d��������e#;��Yኼ���7�H��.���-ي���(����..�Voy��ۇie������=!�A)�h-��<���\��v�k��	V3�
����{p.`*z����m��>�~_�K�q�܃�qT܋a�1�c%��toN���g_���#,5�Q t�XH�I�{��i;����x�O�:����S�l	+e�c$膙�H&�WYCoci��<N�_�p������g|���ʸ��d
G�s�E9�@��K+��(� �K<�&��K�i��J�s���\A��Ey�͒S
jLu�-�	Z���"x��NV�zKTҼh��֧�B���s��+�����*/0����g��X%+H�e��;VG�2ӟO]/��!�b[�XBM$ư�^�U,),��Z`-ׯ��@жm���QҼ���)�)"����x�(TF����1l[m(39���v�P�<����JA�U��r5`ݸ��犾����o60y�-H�H�����m���[E
��|K�5P��@�tXWr2��h�2�A�!�?�NO�Ӫ0�P
G~25����e�te�m�At���f��P�f�����J��n�|�Q�z�����]���yJ�.��0��;�!�~d����v;Fn��>b�M�2�[AWB�K�P ][�%Q��J���z�׽��&����yւ�5�8m�^�]����@${�,���)� ������+���$��� ^H�/��� *̚���e��i:����Xz�j}̙��ǌ;b砡�����Z3�v�{�/���+!o�H7�������i�_�$���=K��ۥF��*o�&(�r{�����2�<(ڧ�>�x+�h3���c1���@x�81�1/��ɂ����R&z�{%x�f~�2M\TC��{v�&T�'�^��,�*��,ϼ��w���A;X�ڧaAf���+�/� ���������,��
ꂍ���a
�r*�{���͢�v��5��^5���$V���x4�f^�1X��u9V��>{��")s}��	��V��*~�L�7\�P�c�a�G���e��0�j�5�=��iK�AS�!v��Qs ��=�T�4�0P9���h���w'��#����>�?d�S��T��/�s���F4dԑCύ)��ؼ1t]BO)�Wm���xT�e��J������Ⓥ.Q�|�\%yU�X(a|L#��J�r1�6�]�F{���!�G��]$;�5pz��;��e�ݢa�)͍'#ӎ�R��É�͕*�(�AE�E�f�4I+b���w�J4+�j��s��`*�0��afq5i>���΂�P$W�
x nQ��C%��=�����3%�'��B
�T U6X�ϵDq:pk�N��J�ZV�V���v�@�}H���:J��M���*�S����w�� �F�"�A
�ռ8��L%Z���u8ƫ���W�U�AL��j7�����;δ�"	G�T���Q��W(���^̤��O
>��G���(��A�Qk��g�4�r6t�g�WJ�5�v�wzY�C��E.�2�Jj�+�kdL�EN���gyݦ��ٺ�8��18���v᷐|�WJ���m ���4v���t�G�U�=��/&I�ZϞ;����lYrlx�.�%pE����p�뽻X�HЧ�2�?^ wWZ��o�ΰΡպ��3!(��Y�(��Yl���'i�79�9m1h��t!Y�g�.�ř��x���Cj6v�'�ys�Q�� �ZVjrA%=��BP�D�'i,��ǻӛG,�N�=���B�l�خ�f:C��\԰}%�txăyF�*5(+	m�,��B�Xʯ�:f\���Jձ&���M�M|��Ͽ�����P�v´/�-6�/Aw�����+h�h��o&��%.x���O�?�n����f�����k���E�g��f����� ۴�M��d3��VU�<{P4k�eB�B ˣm�R�Xo-�"�jh@)A`-�Ļ�:�w[KE�#|�CF��=?���ݧ��e��Ȩ�Q���=�(���aX�"�@_��ߖ�΋P�[G�bc�u�F����$�D6Q��0h*�����g�I�"��GUN���gCm[)C�2\DyA��Հ� /�����Cҋ��o�ǡ�CŤ�	�P!/q�"�k��GE���X@/�Y�RT֗'f�b������o�]��=~" c�j��M-��\��+X���K���f̔ĩ�7Y���D�����2��|!���㡂hzS��]Zf��F�8Qx�̉��"B�]CX7��
�����lj������;��f�'��{��I���>G�ʪ��(�79qM���(w��+��w���s������\l}�}�6���ɑi`K^��9p׿cF���y��w�Ń�CCLO/ئ���~�
��C%X�^�~6sX&�u3#����Q%eD�F/o�2 � dd�Q��  }Y	���WΛd�ʉm�8�|��@�~P�'��ue��ܸ���}��dh�8Kǃ��d�]����?�2�$�P� ���"�ͳHF@�Z�F�����!IA��&�ƣ�Iuȡ����\��sC6������2��B3B�đی��٩G���j^+v'�Ҽ���Ԁjx��b�W�'�-k&����D�<�a�G��Z/j\�Wjѫ	��"�}��s�+q����UV	K���22�>-���CIT��/	/A��v4s��T�@���XB��Ma�n���Ț3�\�^��K�sb:d���'�fY��_��J����\�S�D�~7u;ꔻ�x�	E��Xez��|�
B-Z����̶�[��7����M��X�����q|i�z�!���N��VѭCA����JO�s&�L<�@�,N'��u@�|��t)X�uh��c�CH�u 
z�31G�s��׆�;���	kY�Q����FҎL@ɀ��3���eϖ�K~Wk�]���Z�P����H��(C���_��=uy�"��{@S|�^����ָ�;����ٵ�%ٿ����`{ָ�L쬞M���Ծg���<�V �R�,B5��'���
�L	b6
�l�H]s�=,�B1UEؽ ��o:�C�r�,�Xl��$)Q��c������fɠ � 7K����� ܱ�R��t�pcq?�i��mOϵ.���h�d��
��ȕ�9��T}�˼����@,pU"���8�|=�9<�=��$�;���c�K붷_��\��+eg� 
��v�6�w�4����:^��VA��s��&�� �z���1��/fo���L˔g����(P�ϋ��ʜ���y��t�9hʉ�|]ȕV�%���g�I���osl�܋$���݊խE�3�-}֍.��e�;���?']���^�M����Y
&��(M��^�����@�aG��J��� ���YMA:��O��H7���x�R�M2�rR�@�֩! �x��^�7��Z�>���sj|v���[5.|�I�]���y���,��N�0�\��4P�@X-���d/Z�J��J�q��t�K�	�z���.3���φ&u���{����c�3�����j�����䉆�Ao��K`�c �w ,�x����Gr�x�ƻG�1}�-D�C�3${��n�-;�7�5T�+/�D�J)� h�Y�i���eZ�&�C���N��K��J[֭�X>��F��y/���q*ӿ��X�X5eZ۱�s�SM����T�뽩IO9�*�.Do�oD~��]�c��\_��F��&��ۗ��1yЗ�,�c����0��>��/nl;�LS�x8�����o�ϙ�k�-{@�7�Y�d��c]�<��`��� ztg� ���@L
b1(m�ֳ�G��%�a��n2��Q,��$�擭��*�.��������C�1q��&XqLٴ��/re���]̰��8��,�+���RJ�빲�Ⱥk@��pl0�E��M�[h��i��SɕE(;��C�����?T$z�a$�Z�k���;��P�1�Ą���i>�+�*�Aa/��%L?ѹ�<�9�J�#��RŒ@� �VA���ٔeSݴE�ME�=r	$��W;_�2�rYs�@?��rKoH&Sjr��TL�,�D|�"���7�oa��?xو��@�/k}N���vב\a�pL�T���̱�Z|�`LO�y���<����/>ڛ�&���I����X_�ē����s�qdh��=di$]������-��Im�w��#�H�tBV����!2����(�d��� �/l����c=J.k�x��o?��e��]֙��wF�t�c���	��j5	���hEz�b<�K���'���
q0�S�o�����CJ@�~����&3�}���vy��BG����߂�26T"�@�q��9l���+��3�z#a+gk�}b�f��T}]+�sU�B�9�4�9�0�E�<V<��w��ݍ0�'�/B�2�㌛7U�
!p��VJ�T��6��ԍni�P�>���3�&0��!�#0x7 ��b�kC�U?�HoZs�֒�nY9|͸�L����\�"-h��1�j[A���T\���qC�s�	�M߻�]�|�ꓻ� �7�5�S��<�38�d�o��}וܪ�`c9��:j^v�Z�������侘��C�7�F`� K3��;��v���o۲e�=�uҔ�a�����us�K[� ����N��XR�k5(���h>������R��o���\� ?�H����]fn���ȡ7%4`L�Wz�u.�Cۛ��'�Kfm��mO'�%3M�˃C��T�����U�� 0Z��G�>����=�����^��,���h���d�G�lP�Z�� R�R5�F8y��V��H�X�� C~��d�Թ@���B^~!X���Z���_��9?݆���ܹ~ٷ8�����MREt��_N�A���Q%�H�����:�V~P�;��S�,��iS�b���3�?@�2���nܦ�T��J喑5Y�`;���j��̖$[�3�5�	`1�(d��"X6�PԷ��]w����:��4�Y��^n.�a�	R`�b�D��5���	�s���s{E��~�5�EX�*��NX�%<'�?��Z�qy�s1�+ȣ`�F����x�@Ò��d��������'��lc8&P�X!�p\�5�놦��嵍W�䗽�m��A���eM�73�:�/,�N5�/m	�;��H_���*��ZJ��� Q\#�&��b����^����J���*>�,������i�A_UP�FX��6��\Xe)o�7)�F�a��R*դ/b�[Ba�gӀ�n2�����,kh����F�M)����q��u�6R��@���%�r�0Vd�xJ�%ޏ�<:Jp��ӄ\�@��j�����\r�GO�B�$�Wޑ�q)4<������|v�2X�a�`�pۮX|���4h"1)��0-�:��=mq��ƺ5���i�mB�b@�7����e; �:�w��G��%2�}��p���
.Q��~'�G)�SD�@{�Mg�)������˚{�E(�4��X�[�Bc)�E 1�/�X�O�W��ǳeT����~h��o^�	с��l:z�I��6=b�J��ZN���gk�8tXc]��I� �(T6*�Q1�Ԛ�{��`����W��AC��,�]��C#�ZS�ϜbҦt�� q[���ϋ�L*� � 0g�g���c�� �VoBǇgYVִu���L���f���0�<"��a��Z?%�	�:��k���'��l���kp<�k���5�½3�q��,�)���4��k>�Z�\���V=?��V�� ��4O�Ǵc�`ԯ�M�U	L�������]0+ד��V�ݳ��*Uq
��]Ore�����u���_��O��w+�~��Ȋ���}��ٵ��5�|Z�x9�����d����(�[�fN�)?��Q�-��2�إ$ݾ�Y���Р�����ǽO�7-;�����Ġ���q�
>i��4�S<�� �����L���X>��K�wr�m���yg%�k�7VD�U��gV�z#�g	�����Vs8Z8�u��?��X���գ'B����k����'i��g9�=?�J�6yu�^N�)���:R�Q���A$#j䂄1o�%`�h��U�|ī����Ϳ�GX!�!{��*|��D-�`�l�</��#]>���,��z�K�{|�����D ���I7��� ���C5=������Uk�3c%v>�MA��I�y��h+�����~ן��%lC�qܫ|�`_�Bd[�vϞ�o��'O.2�'ܒ�z���K�A����v��Pj%TB��9�IQF����ò����L�ν
֭pU@�FT������.�����f���Ԝ	�.Q��=3O�X.����/�CM�M9��C�}�jh�O�el��c?�$M20�d�s����G}���?:z������@�`L=�^m�d����V�yRxafA��j7�0���r�P͍s�3���|��/���]z6ޅ#뢆�އ��@>�d�Ye;b��4�^����?��м�lBڅuּ߯BzEEl2�����a�qC�� ��\��36����4ҭߞ�����G>��.�{�H�����1u�t�g�W� �y8����tL�WԽ[�%9��}���T�y�[�{�EBq~���R_�
Zp�ռ�2��;u���TF��2uѬq��G���%�ɽ��_�wiz�d�p�����,H��N�f#y�'s������[,}�.#2p-F����l���ǥ��$�妀�,��]YO����j�e�Y��a���*�7ɣ)A���&~B�2)��1<��b8<�m;:iץHu*�"JwȠw^�v|������v���$	+��dI*O;��:��3�U�����Rˎ�֔s87@�ϟ�O����q&`�\̜�- ���ak�Dѿd-��g7q��)��aSdjF�\./`���G��K��٦��Zm~����Ù�>'���B��E�"���5��G����$����F`�O���~���0S�q���5�}�ɚ�O]T�s�DʈP����)+u�q��M�/�9��#�����3E���_�Ru����v�� !��J��Ii�o��9aʅ���X.8�� T�PK"dX�e����}��?_��ߕ��ɑA?��D�5����	�p�b�B��m�@z��2)�a�N}r����D�c� �aR/�	W�cx�$�j9��		h�������
�߶�=W�y������rQ/��ԡLrJ�cR���.�D:�Y�'C�⠖Co���M1t�X6����#��j�d]��o��sKԉj	�B�s�]@�NY��(�34@B%�c���*F?LXoW�_�/�)�҉���k]�"�*��XnEf�D�y���5��hv��RDȚ�$`��)��[�UMAT�+�L�������
�*G*X%"��n�;ڿ74�-��y���oq�D?�."+��M6$J{�ܣu�`��z�0yZ��(�u�$?�{�K����D�胐5��a�m�)��+���S��%�|���]���ږ���t�+6�s����+��9�a� �b���q����a5[�w�7��Aǈ��ǅ$��y7^/��*��G���}�BY�D�>d-���=3͊�;��J����9ȠӁ	_ �``�>��O�d_�B-K�:<f�yղ��o��
�x}�;A�u�^9�(SvW��w@g�&5>�8l�z�n]��}4�l
rߺM���=��bJ����Dk�d�e���9�/��\>�eE+_�3��;q~8Ov�4�Z�D{
�� ^y7�',A�cN��������O$���"��;-}t�˰
ڿ��t� -;#���NAMa�����a��	ȍz�U ٨�O[,+�iM5V��t�,�u��076t;�>�rr��J��fM%�K�hr}ߏa��� �'B�D[��B�P�V����*�н�ȍO�.b��TO%m����-c韱���o��-����	������6x��m3,�&x�p���5E�P.�b���e�㶄��6�!��iz��^�1�Ɉ�bS",>���З�k���2X;�C�W#Q��-l�:���i��O=�B���]s=[��ژ�_��!�:+5��<�DU��C�s�#'��
8�X��	�Bc�鷃T�D��(3����.�0��ô�T�r�VV���װ����G�:gT��^:�����u�A\���Z�K�]2���u�Z՛!��4�`��\ � m"��xMs#�ۆ��HN[���;�jJWZ3���ށ��E��q���� Ů��zk�TAQ�4s�#��.E#k�A�+��0K?� }#ۈkJq���l����U{\�`%
%�~��8"s�	�ߥ`җ���Щ��rY�G8��̳;[��Y����gP4`��ry?n��}u�/�H����"p�Q�<���a�쁡���}B��T�]�u���	r@�
`~y3�Oٿz��ʥt�ҥ�Xv�9�����!�+,ݏ���\�=ga�����(Ńx����C[�k�W��������+����q�i�|��xt� U��I��	��M��nO��^#H��Q��9 �sa��lQ�cCI?5�:�r��Y��7M���m�BV�5��&a����4���LҰ��Tx�>N�;��6<H'�*�6���sN���
9o�_?h�U%���"a�~�̓�f��E�A�p�ZI���
�á��2�I���w^iO���L~�ޤ�"�� 5�����`�]��}j��`Q�\�����X���?�ۄ�P1���{�� _���U ��|ո�w�F �����V!SLo���Q[A�]f�c��)\5��Й�&8��0���e�)6f�٠
��~L�>� ��<Ջ����:\��2\kڢ�l?	�26������D:�(��d�a�l�yi@�����XԘ�w�ji���u�$��:A�3�!����K���k�뮱AV���!(��'��r���J.0vwE7�+�w�����������`��3�_�����_�� �E�Q��J5wG�i�-�E�5A����;E	n��Se�Y�Gܠ>�@�N�RK%F��!�<E���щ���-Rt�x�C���$�챶pՉH�Y�]b[v��fw�Gw�����iI q��1|�6N]�M�+�cV���+��њi�Ư>4kzP%A\QL�B|�-��;Sb�`��T�-�Y�����)y�v 0� {�H����,2
x� �}��uKK���*��� �FG���IY5I�8vop�ؽg�hrͷ6Z!����Fa�Nq�Y� ���"��;���'$����"�|��E�H��D�o�̏8��ej ����G��ZyvDT��Pڭ�|�=�$�K.K^��c�.��=P��$N>�O,-�!�c�$���P� U��0c5f�|��tҀ�����WV����s��Qr��$B�3Y*Q;�{g�~�$��4�k�-���v�Шa�,e��Y���-)q0��p���
�JzJIc��Jʎ��TDq��=����p�Ykq�o=�)O�eнǧ
���k��y]V�Z�U�;rF&)�-?�T�F�N��:d�&�����q}�w&Т����YҔ��4�&��Q�0������6ožC��\DH�kvS���O�
��4u�dC��
�P�J��V���%�̠2�K��'ź�@�#�WYʚ�X��T��`���龲�<$�4�Q��>+�����܈�OLUi0/������S�M�;T������Ԅ���2]6ٓ1�%���*
��%��r��%0t�7� U@�j�N��V��e@�3%Y�1ĳ]�rb���6�b����v�c_�s�b��'��6v�	����k��ws<bD�B�v%EM �E+\�SшY�;��-7g�48W����y�Ƶ"��*]��|KUa�^W�6�,�׉�K�#�Jt��,����/R�W�f:��Bq_���ԛ�I��m�%�����*3P��\���PE���</��w�t�K����K�o�r���-\�b�I���������(�L=l4�O�M�u�NP�F�K"+���:�^},���x��6ʉ~U�غ&�=���1��!M�G�	�W|���2�e���ts��m���9�.}����
,jk�+�u)�)Ȳ��#��t��m^�vHo� �9uE�a�ݹu���3B~h�gY�Q;�5��D�+��(�F�HV_k�:��P�� T�a�h�|-mыi�?�v�M�ި�k���[u՚ҵԕf�
��lt�W��-}�>|ǳӊĔ�M{�|�k�d���Plw��M����F��%b��O�g4��
���Z�=H@�|�Z^^K�*�i��N�4B�)����m8�k1��d贁1�X�����ȼ�L�WT^B�!j���ew����S,�L�)m�@�O6���5��I-)ko.���u5��H@)���/u�M�h�{��	��;|�}��W���d�V�_ȥU�s.4�:����<�'qy�j���D#��c��b��n!x�j�]�o�W��YS�l�j}`��)�lnE\E�L��jt���vKmT�h/t�1��9Yݤ��x��1��]�`i�D̈�/(Jy�t7�vb�6^�����$�N%���Ri�Wc�+y��ek.���"e��AW��ĸp�Y|�x,?ᩋtR[�72���o��b������It�4��a��&:�z�q��j{&�r^����%S���_�=�\�vk�s��3��� {A�Ί��Og��,����ʿt���o	= K9�u�Rv?�>�ۋJ�~�WJvS���83�3wy�|/,�o@
z�V$ʣh!�z'�408C,Q�����tn8Ͽ��4
oEz�����}b-��-�A�Z����\�0����o�B����Ⱦ����wm�d�|Х��#�,����+�O��K ���r�u1=���c|�}]�ܫ��:���S����;xu�rj�QIZ-�k1�1�^ 8+�v2"�ʶ}�0� ,�2:�f�G#&��
АPJ�FL�gw��r8i6�j��׿��34)���j����G<��N�·$�lǏ��w����ڛ�m�g>__��E`��z�+�c�a��t�Ҿ�ϔSG!~���	��
'#��uÕ�˵��)N�,�'A>�Z_y�/m,m�Š�{�C�E[�sV��������Y��{P�-ڴ�t�gpz�P���������&W���O2K�9ڣi�E��EC�6��X�M3I�ԙ�O�$ۆL�'��,�;SgţI->n�:��G���y(��[T<�"9E�4����'�n��5�2{��� �n���{W`��F2FU��ܫ�<�m~�[ b��E#��2��Dju��c�'f�}Ԣ��ce�܇l�uD
6�xK�.�"�guQ�"#��2�SQY�c�n��t�ƙ��#�mW���o�ێ;{>/�L�����Oe**��Ǐ��[�d��ix�����Ͱ��_y��be���檬{Z�l}��(����KzZ�[�� ���'װozT���"��^�*eU��E�����\���:pm����;�#1�ag�d6�Sp0O	��ͭ~�c��1Ƒ�xx����{��ױ!A8�R7h�̜0:v��o����^N�,�R�����ރ3��'���Umy�K�| �[T�<F�qlY�PUVdV=Kk�� �+���!�~��D.�h5C���y��8�iU�_�M:�{�_R���L2����UAU����.P3Ԩ?����KU4�=��4;!ĕ�X����J��
Vp�K\݂Yei�/�����2��2�Tc�p,�]K���/ȥ�F�7��y���U�:�=�j�$u/�1W*��v^�l�����3z׫ w��V]h|}�7�e�k���)�	Hӭ��~'�}��$�: �i�,�r�D��D����S���ֻY}�w��ᙲH2=�X��o�9X��f��g�g����4�Q�;)���o]���Åxw)5��K b:r{>��ۍ��:O">���*��x���~`<�-��?��E�b���ӕ����*�J<�!Te(.�{;=�H�h�ꅷn~H��O��]J�²i�|7b��@}[wy��.�ñ�ƥYͯV�W۸H��C�/�7��S��|��;��5����,�؄۽��h=�Ƶ�o�L�4>{�Q�z�����`��(4�ⵁ.�ȬK��F��X�7�����(�J�5�7݊{�G�+�����3��CƟ_�	��H�n\s<��� 
�A����|k!���A��ƿm;�E&=�,�
�ݗ�󩂶BF��/�@�C:g@�aa�:�����7��B]��
K����$����_<r�D��M�*�;��W5�ی�4�譤�����8�d�d��|�mc�j�M���L��	�/an<_����:���(m�1�*��8=�5;cw�@V ַ�߸����~��.P�0V!q�7h���q��$���\�k�Itn/I�o��"�ӳ���wƈێ4��L#I��M�q���Vӯ&<5
���"P��Z�]�v���zmp�?��F�POd,b�wu�y�tr%K?%\p����]8O>u]�-~c�nǘ�z���S�<��Ws?6��r��+�|�ĨB�ˢ����>Y|\H0��7�>�"�>�K�N�Rl�u��n'~QxԪ^�"С�����	i���Q!����3(�-D���.;Y�ԣ��������;m�.�43\�63)%Q�٪��ϙ�Xy�����������)D���XZ5<:��L�W\�ι�Ζ��C�徝�B&(~��)�(uM��B�h��e���y�g�k��<Wh���!��#��U�sGY���Zn��&��b�3l�Z���a �����P��P-�8r������=37H��.�V�V��a�`���5����n�0�{��/�P�	��{C�T�_{�}�Zޗ0��ܜ��8�K� �U-��m�����h�����U�`^�\	R�0)V!�(a'��;�+��n2>f�X"2֖c�zL2���UZ]�$����O���
��l�A��֯�߽���#hq�x�@�4�ت��e[�DKrv*���wC���Ha���S,�ϳ�^� (�������6��P*!����}<Q�'�^�I���m�*D�r�#d�G��i�iU( ?`���!X�I�Ԋ�����~:�G3�Ц�x.�(�
p^���8C:�A���?�84��&��<��2^�+���:�8�>㘻��a�o���<3��|y���8v�,�p�Ɠ'�����8|ISia�dr�<���s�]��ji$Avh��ל�E
x������w9�����1����`@9���O��~$���� �p'S� �0�oZ��s}�J
Iu(A��tݙ/C"H�͋�h׋�4���樲�X�`�V��>{�$0uEa��3GdE>Ғ�+�E�B����]o��P!�nxp�����Z������Ô��?�5+t)ӓNH��I�@�]ْ%��=_z���*�`��eC؁s�}��ɑ����� ؛��\e��<�Ӕ������ԑJ�?���IC�ȧf����K7�,����R}�e�u����
�f�X?�e�Y����]c�6q���uż"��|�𺸶l�i1�'d�JJ���-i��q�X��9�9hL5i�h��Pb	���h+7�� ����C�!��:{T|Ael��`UW��F@p�X�o��Q��6�@t����v������џ���«��T|poE͆`!��Q\u����%��l�vU-��{��a���
|��X���Q�h6�*��
%gLK���sZ+�;�'Z�"����J��Z44+ꋛ��<��*�TQ���ϳ��G;�v`r����lF� �۲��1���T�\��·K�d��psQ�%`�r(����s2e��EX�>�7T��ra������.u��+�eud%��蹐�9K[�z�ik���>�ݓq��f�����p�,�i�q @p�B�90CJ6?���J2'@���f� �u�mk�ւ�6���ٙ���@Q�>���]�n�n�.#�m~�+�oHJ;� �|#e)IN��)9��Og9���6�_K�_q�Y0�q�r�[�/v<��YUH��	!~k��"(�rl�ę��� ���e�_7���%�$�Ψ�{�2������iMV�ke�0=t�@�[z)'�Y�NC�ݒ�p�ͼ���/'o��?�{�x��Mu�y{���$���s� �&	�I����`���Y�j�����	��5�>�xm�+z�X���9��m���r�2���*],H���
�1K�c��h�wI�!�`��:�B���	�#mǑY�͓;e[�ܥEи�ll���{��Ο�2���>�L�t��S�n����n�Kj�XX��� j─0�u���2�K:�s#]�;:b��e�eaQ>T��P�BqL҇��-�Z>T��";ҟh���y�ъk�+��[��:P���I����"������yI��X4�^s���4�d>�(L;^�߻����"~w����(t1�u�%�R\����E���vq�O�a6�K?�*�t���Q���e�ȍ��k��+DVS��6��G�N�O�"��i�ٿ�+�����4�1��uȦr?}�&��9|;����t��9R6F�YJ�� i��.�i��[�rj�D
 {�p�j[�݅�v/o"�E���	�o)` �l�W#�P�g���}z�	:?&���,N	n�` c^F';L*��OLVlȆ�T���܇�Fz`/C7j1!�s���� ��]X�!����G���ͯ�ZP/E���Z���\���gs��m��=L�
�g�G�.j��]����@�8�(L~s@ l��vzJ0����)�F�7ECz��HB���z�6���f%��}�V/�B��W��na�>��OV���28ž�	t���"�v�M*�xϠ}߄T��A�b~�5p�J��\(,�o�����G�L{���`�˺;Gڗ�B�J1�������i>�Ҩ��	ED���ܱ�(�V�G%C-]��>�k@q7�ֳ�!ˑ%ԁ ��R��ADp��R�H���g؊��б�ga	]%�k����7 ��^�ז� ����#5��F����]�n	������< �j+���;��ֿr�+���L��N����������,I V�lni��m?ޢ�Q��]��;7>����*x��\�E�y1衬��bAEu,D����'N�6Vv$�";���!�(ȗ�NS����V.��w�{N���a>�5E��.Y�EB�+���V��=��#��R�$g�s���I��~YE	�ה���
"�"Ǉ�e�H��{����9~�2ER\@{w<.�sCs��l���%�w"��l�,�/�=�W0�D�Ó<*�j-���&�XJ\�o%��}����jDt+~֢c<3���+b��4P�A���A�#�W�5�j�V��_��R�l�?�;�J���'��S7��g�\:}1���Ab��Rg=i�G�[���ɶ��#1�[�g�����doY�6ʢ-ϩ6C=����zuHR<pv��^�u�+���u�E��tC;���Z�i��T��_�\�U�B����iI
��J&.� e�n�#~ī�}����D�z��+�!��Y	q6X���#O\��y1#��Ҭu8;N�`�g[O\�K����z���uq^6�u+�=ㇳ�Ί
�	�����{���P]�BL�+q�"�!��h��� ��h2�y�X�?Ym��jVU' ����uY޼5M����^�׈����Wr��H�[V��4�iGFs��8�����n�Ր�!RDZqoj��i��Cl,���hX:u{+�B[ɍ0뿱����}�S�����l���T�f/��Q�� 	k��>o^hx���
���$�aL�Ul�GN�	���y�����QduB�Ո�K��u�g��B��O�G0�����*HP}�o���uU�Rd7.$]H��}�F�S��4��k+�Y$W,(8��X�5�� ���ߴGQ�����rls����)�~��SXmI�~���~Nxo8ˏ�`�� Կ2�r�?��;Ŀ���m��ȱ�w��`�����'[�9��rY!�;yzr+���wW8��[�{)��n�8�z%W#�RWk���.>��C��蛱d�C%gF0>!��kHE�QΟ5�=�5��{��>���ʥS���s��;<��S�C|:�,���>˾���܆�=c�l��<B����P���	|�B�ڰ���!S�A�H��N?JV<�$��;��*�6G�����}�wh8�{�E�0��/�T1����������O��MG��*�0�lM5���h�V����%�$�:eròp�C�+�|��$�Bޅ���H6�2*�N�	8�n�#����"��P��B�r ��S�-�̊@6��E�	j+�s �~�D���V��4������op!���7�"ސ�z�wPZ5Mʨ%	�S��]�\���y$]����h��E�h-#����A��o�@�ʬ�ŏ��?��|��cE�yzy�ڳi����
K���^2UxLy���hA۟	��58�ě��I@��z/�k"	��)�;0A�pغ��D��N\�	/��XL-�+�)'N��HS�pŇ$Ce .>?���e�]fy�)M���>.��10�ɀ�L6���喂����T���Òzu��b�9~�J���r���R�*���
���x�2�nɡ/o㙿�'���3^b5�F��f1��/px<����,�֕�.(�!y�������+��Be���Ck�[�a�k�� �A2~�vz�Tn�� ���f_�:I�2;�Fy���㶎F{�&{������KVDmy���oy�� (�O�bB�_�5��Z�CH.�6�Jl�$=��o��:0#d8��	xz�w��2d�"�ӹ`�6�g�Z$yj]̡T�H�/�4��7��4_uZ\�47����Y��QC1wJ]
��Ɉ�"�Z�������N���2���"X)�g���	O�Q-�3u�wp��dȠ;��vH�5�y���_B����y��%�_��<�8�xA����GzH"bՎ~�Oj��͹�5�tn����lmz�,a��q�ى�\�L�#W˙�BE�g>&���a�1���Ӗ���3#V@S~ߚ�W���8Y��%3�sf�(��6�pD��NQ|O�J�p#b�,�)�N��瞝7�bٲ�|�Q5T��K#yW~5N���G�K�r��\PR�����a<xJL�악|B>�E���Vj�^w�������N��O�����n]�1!��:���9�c�{�>��X�`�Q@�6��M�ƪUM#��Hc�".ZG���nm�:�ܗ�]��(O����������g�{n���,����K�&ч��T0�����+%�u�Vx:~ ��>d�Ȑ\���k|�6��������]����|��r�]R��]/ׇ����%�.4��B\�`��[�e��d�GáH���&��ż��X�h��q\��D��&����+;Jf�Ph�4n<|1�Q����(}��U�U��_h����IW��W[g�͚��m %kߏ�juK^7�`m�
��NE]�(T���9�A{ɽ���n��e�WB}��9H�#Ai��<�&Te��5}�t{ځ� yA��������h��Z d��t��[
���>\/�%����s�����&���e�0�Wޓ��4K�h�� ���T�Hә(b<*Qйd^��$�~/�����)�؊��r̓�H�9-�&1�Δ8�� ��\�JrBb���sָ���-�v����M�T=ߥ}�h�^[�s���Ⱦ�/�Ƌ",�T�����]���(�ӊ�T��5�>�� ��_^ax,C�(��i����^��Xw �E^��K�7[�ӍCH���k�ʴx�Z�����B1������cnk������"LW!���C�o��.Dq���I�G�)�b+	\kF����|o��*��s��"55b��������^2` Y���p�g�����a�ZR�E�:�I׭��Y�Ͳ7��[m�����(����*�9���Xj��<�>m�g�P4}K)��o���z��ܢb2��z����ƹ���g�n5�FhBu�k���=��6�M`�W�R�3KŠm��&�~} �Ǜ�7�}�b7�A#�J�h��|�O9)=����3�#�߄D�0
P��R|T�8��di��+i�h�v�J��9�?��sw�,䑼k��K(�1�-ɏ�� Q��=n7���l׻�	�i�1��A�xT^�ֳ��Lf���걁2�W�!�%�2`�-�F����m���T��?�,�� �U�$�k�!.r��7ܽK%��4Kx�)��`󁾕R�b�<<A�lB�l��5waӇ��?ꏢ�]u������w}al�N D�QTU?*�7.�{�єٌ�Q��vzj{�-hvmw�����t���:����%�ِ��퉂�V5��(9Z;��RZ����R��}ho 
��z���ޖMI� #�S�_��Or���6����IT��Re�C����T��a�ӥ�\."��~��Jc�'��>'��+�X�^^�)�����|�����|��N�����>�|m@�o+��#�m��B%�)�u���,x��t6�����f�W_8uvK���ݳ�:7�o�}	�����cj/��3z�i&�����ydq�d�g/\�c��w;#G�4*6n̉�}<A��F��+;@�̤�3 �f)�ݸ�v����Hƚz�9�%:��_1�or۷	2������Q΍/*L$B(���Ѓl�@�u�[ROU��8t�(<��ç����ċ
�)��Խ����U����2��^�񣍆�9�QY��)�K��Ú6q=`AM���\�F_�H������ހ��\�K�>��L���@�0T`�ՙo��T��O����`$A�"� 
��:B�����3�؅!�YV'ɥ%�v�-��߭�#DZ[6� �nVD1
��`���HI��ЂJS!�g�W��e�����<�!�5#�z�
����B�Y��_�\��+0��S$N�(���/wK�� ��Bҥ_�p5ZI��[c���]hA�q7L��^�Ԇ�jűC��O���'��6�\��bI{3�g�f�ޗ�Yõ\�'���d��6�V*��Ӷ��tVk�Qp�su�BM 4,w�Z��1�u�3~�[���+㘋cA��ڶ|�Y��,���g�J�o�.!�&`_Y�匵pcbt�"�x��Q�*�x&�Be�K���3L�&�(j(����ȥo?�L���Pc�XE'v<^V��q�R���0�'~�]=Z䞕/+���i����].1��Ri~r��K��ź��(Ķ��Z:�#���XY��(*~��n��
3<�A5�;#m������3�
d���^��{'l^��1��v�5]V�Zd5�taM`���MxضIo#�pŮ&��;�e�����t�q�B��q��
��=+�8f��]�0����)�����t9tǎ��r}�R5w0ZZ�@���	*n��	���EX�f3w��@���5�%���fkb(�i�cH��ENd�˦{��~[\��2����R�M�#+��oxpr��~	1st���]�~�It@#I���*�� �U�3����_�rA�R�v��pͥ��Pu��\��|sbiv���D���}97�+�f���*Ť��Ϣqsx�h��D&F���$p�u�_�g<^����+0��m��)�$�a��0;�����nay�c"$݆������5-�p�m�yF�r��ՙ�
�1\�Z`0N�/���N��k@�'�U���Z� *ʝ�PZ�� ����٭�߭xPu���i�h�O�Q�%���C^�f��z�\;��
΂���]P/v�ɏL�T��	�~P) �J�^����)Sd�| �H����dwȚZ��=m-�����9
k�w6�p�)�w����m������+T�`���T�1�Z��Hu�p.W֚�)*�Cw����O�(��[{N����N"��{Zݻ@���la\���R�m\��qM  ��鰯	1���vU�Z���3:�/iSW�¾{h^>���F("��oi�u%+d�S�����"���-uwAG�cn4�E�ܚA`�
d�'L�0鴹����0��������U$&3���j�����Zt&��c3T�!=�%��
�i
��������pȸ���Vk���"�E���J�K�q�����:�.j&I�*u�4�ьm&�x�zY��#��i��j�A�����l�-��(�x�
��>��
=�@E��
����g!�{�%�]:��+�q��g��M��,}sL�A��2�À�1��dc�>�m��O]
���穘���5�&��c�R~�ա����3���D�|=z��i�˄4O?��8zu���N w�������+$}��5%�t^i*9�#�#�]Y�\���֗7a���փ�A1w�\ �&�f��L�`a�>��#�i�=,�y"&��N���`!���}�@�X�Ѥ�!��;�Z� �:��N n��	��4�H��u*�t&���]-�o�3�Ɓ�ϕ3��M0n��#�*(S���u��:�jl��R�����fݡtA���ck��0!�͟�8^���tߑ=@���^R������)K���)UW��2[�< Ѐ��Y����G.t�䠷S�0�H�.f�I��zpY�����jT��4���I�O�~��4MQ���`j���M���� XK,njrqz!��@iN�k����5���`����?LXq�&�G=$7|��N�[�}IG{��[я�������b�����Ld�C������zL�9��٢��oR8+E1��;ߣu[*O$�#��S�5�Q�J�Mi5�i�����}V��n��k�G�I�h�p�~�-?�)5���������:�"B�Wײ>6zd@"��C2;�ӥ,�$��^�MJ0��.HZч *O;-�~|y��.������Un/y=s��}b�����
Y?������8g)����?���l2���q��Z�e0"Ȫ��J%$7W��-.�\)�l7��� ����B1j���l�A�ح��\�lJ�Hd�25���z$�@��燂�M�j�L��S�
�g[�-�̬�~ϱA-�!�����&\eZOaoEdf�?�� �kf'����MWV�r�O�[��>��x��@ԣj�q:lBT�f}i�"��{Gj!$",dALh���R�k���Y��g����5�E�����������$����n�Ν%v{����������"�9�h��q�և��p�u-����B�AJ=��_���4�:�����W�C[\��d�w27Nt��{A��Ο.�ִ�������3�M�B�@���a"��?���į'�,��m���KE�G�3)WohdQ�`u�G	�w��J����p1�H|DN3v/zf�BV��#�|��dU���ov��*��@����G�s�V��6SЖ��ϻ���֚�R�P)9�(c�"g�<+GflPB">2o���|�Q0�~��g�_v^cKJ`�oOJ�IN�(_�O��3�*�"���6�ļ�F}I ���T��u���Ä[�B#�g͵7��7W���kT8#���j�h�oR.b]ו$v���`
���Kv�sg�Ui�6�L@���b�.�n��'T��z:��}n�Aǔ3L��k�`���b���[B�;�ǟ����;
���n	�4*[0A���Z=đ^r�?�U!I;Q%��2VQ!�	���K��2���ݫ�sP=g>�D(������|,�ڢ�!��D�s��hE��h��CU�/���q�(F>���>���ć��j�:�������ؾzC�/(YJ)���,8�m ����IO+4^Ki��6:��n�5�.	��� F��WY]��	
�q{"��$���J#�v���3�����"���FA��8��K<���'�\����] )��Qm�*6� t��ڦ��W���:?�?i��8b���2���,�C[�0���%m?�zAnO���u�s_=P�㓚�Q���T�pFG%��E�ZѠL��2�
剃8R���: ��x�XI��lb�օe4p�P����γq��6s�]'����\��H���!.�UAfphs'�]n�q��D�1�WJm��3���}����@��=T������o���3��l�N�V�!q�ykz�>�:p�N4u��*A8����O�u:J�1�ص��
`�[U����Ov��t�4V�I�m<�w�cW�/3�/���a�?N8���J�3�'���Y���$�h����N�sÕ*܌\��%����﮵��S� \|9J���4�z��AU̔x�����OF���=�Z�ar��aV�$T��ܙÌA�4���`k��/����}�<f1;D��>�>)�yiQu�P�]e�Q�(�u����ڋWL^�E�	�J���ԲыV���M]�0��v�]
�p�<����A�y>�p!W�I�ӵ�[�{��xt��xfڢh���s[2�@zK1�U���6��4Kf�D��=C��o�į��ː�(����gxq)�s�>抵���6�Y�[Y?m��P�~t��;����&!*��:w�Y������X����	^���H����кV���1�����R��⁵`��)�y��ѻ:3�78<�+��@B͌�rVm<��f���,PX�-���k�+���x�"��{0�6&XGi���4%G�q�`a��?t!y�őދz��,N��MB=Ez *5S�@����<�e���
�3Y1��uާ����"�z6��z�)�U��6Upd�sJ�/��'����}=,cZ�^.�)�C)�h	΁3-u����h4�TZ�;g��uؤꝱ�h̀8f
M P��!RK�����YR�� C=�_G3tI�qRNz����bA��ObR��~/�nM�xwpg9!���.��6�`ӑAN[��x�o���������6Oވ��~R�g��_Q�9����dG��h�u�{��v��ԋia�R��[�Y o�ܛj��Ӈ���6�&�[a5�䈀n��ߕ!����`y'ۮ�>��].���GJF����3G�+�)����
~<��p���&oP��
ɤ�ٱ���q�1��\�C�_�^�J��a`N�Q��,˚��1F�:3�
��������]ձyI����[
��r�R,%f�0Nϛ#c4pתdu���zo��a9<� (�԰��p�'vv���yX>�#'@#ٳ�>ARsσ��3^� ���Dw���G:�"��/
Z� � �RK��z,��,K��!Z)�-�8��Gu>�MW^� 4��@��ap���?{}"���V��{&��x�H�4��+�
%a��O<kw������Su���^�Kh���RT��+�ÂyT4�|��<�n�Ҝe�[�����[�Oѽ2��o1�;�!����|}Eb���c�����~98 nBf��q�F�� v&o��Ym���Ak�q>�Ӆ�7����B�_p�����n9v�&Hst�!����%���Z�=�7uj+�eb������^^A�T`�+'9�>䨌u2F��+�(��e�A�kX����)k�!�J(+u��O��?�8M�n2���.u� �?93�V��`I�q��4�c�4���N�*��<�~T�'T��'c	
�btf����#r%��п��6u8����"%�&�Q�[K�0� i˓2~7���V��F�G�D'6^8�9��p��)H���t�)�?��E|c�K�gm�)Sz;s��~!��J���B�<�0o6r2��6��-#K���ԺR�m�E��w�\-4/��u�kպm�./��m�E�Kw�D_��ک�JB3�>���e��n�-�	��곟��^��F=��س�)�&zF���Y�L�)�������� �h&kc�{GF��o��g�R.�Y��l�x��O:sk�wd�}�S&�+�q`��3Vju1vg,���9�Ӂ���cb�.�{B:`r��s��!��04rZ6����i��0� �3GUv��!o���~"b�4<Þ��ɤ,l�k虷�>�O�j7�J�
�`�[��7"\^'D��z3����8��s����-�	m�F��*X_�$�K�����D�<� CT��iX�]���`C��S��}L��tT'��O��z��\#\}���!��E�B�����<�Y4߰��q�6<lD��{���ĉ����Ͻxfmtȓ�"�H6����aރ��Ku��!:#�z� T��1!S���o TD
�x���j#;�!3�h=4��I��T�I@й�I=r����h-B�AH�@���|T�a'����Q�#��v�����/.�F����Qą)����ϵņ��?��p�ytB�3L>/�?���(�_mivU}��/���� ���OʇzR�M&�v�����)��hq@ݲ�GJ�y��5e�v��jg:�aR}�^e�	���ҡ����/�n���lu��m��k�Q��|0:�<����켵k�X�3N�s$P�h��(7���� �0��T����)�I��=�?]�����`u��ۧ�uD��^�ӱk�)n����Bn�����9�b��=j��ۖ����ł45f	�ʙm�n@���Ed4v�a�D�����MpX��apK]���Q;$�/��|o܀�2�Ś��<���,qN1�0ʝVgQlaآ@�@�"���G�(G�Ϋ�"+��[1��=w���a�!�X_�Գ�<��G�1yEqEFz����u"-�[��VT���9��85�ͻ@2\��DѦ�(� J9f��'���"�_�2x�N��b>B��qͶ�,/��䱃mz���X�1��!\^����2����#�Uc�V���.-4KR�({j�e��;-�l����RG %N�j���L��%���m3G��|�ΐ��#.*l3¯�f[���a��䉐��{�ُDw�"��=� EL�)z[`�e�k@����ޢ]��Br����l�=4l��I1ua��qq��2�n7/����لё�����J����H�������:1�q�|>Gƶ���oU�l��|Wd���m�]�ѺY͋좳�L�4ԝ��E��_���M��T�P/B6��0�v���^!5&Ԓ�j���@�(Ԉx���? S��?" ��4��mS6X�)N=����pηuR�O������Z58܎�Y��H�V��~�>��$��h�8�FK�E`u�����PS�:�b�<6^;e��.?c�C��&�P�&2�J�.�Q;�?�� ^}���/���6%�L����oxt)*}[z�G��\�R�����|��Y���O2Z3	�Eh�iiw��[Gk]��<��=��'�l�-��?���X/�������|��Ґ_�0�i�ŵl:P<a%��~ʣM�=`WB�i�m˦��Xը!����#��h`���cE���5�Je3�R��zC��I�����x� �tԣ�3�t���>[@�7�dÌ�.C����j�bq��|	�G��oׇ������F Yq��Y_ha`�F�K�����V���1��$�eʚ/˫(����P��pp� b��2P���w�
�92�?�+�!ױ�$ܡJ���EKŮ;������v<��rP�*���3�⌛m��,/>B���w�'0�8l|oQ���r��KS$��Ƣ�Q<�⎕���"F�iy>���������I�dN��2�"�MD�ɰ{���i-��y��ŝ@�`���_Y�
�d*�T�IXx�@�QU���͜��.8!�?$��$�!/9ix�R���=빂\�o�� �-&:�1�u�,��p&�!F
=C�xo{�	���Z}4��Coh�L�8�tFj����Ó�*J������D�H����6��4���[��ն��� �0�v�u�JW�Kl�Vf��Uo�5ϏT�4l[�	��D�c�1���"�� �V��\~s/A;��WC?��i����Vq���5����#�'��!�F�j�2�~w ���9����� w�����3��H��=D�Cv>im�N��L.P�WJ;���Snd �H�G��6�Ej��XL��ZĈ��V]��tj�#��E�%wqe���|KS��>j�|��솉2�;-���rp�!�qh@�Cz��v���̲��L��c&�A�#ź�F��T>QIGtA���o+����	�"j��٪�?g���?C573ַz׺3>�H�l��M�L�Y6p=�]&�L�W�orL��?!�5 q��R�UqF�UU��7��<I0u��U��3P��Y ���<�B̾1�5wA�n�9>m| vu�Bs��&������¡�� ���"�4��T7��Z���uZ"�� �t6y7�R���8.��Ai�>��f�^��lg�vGx'+�X�v{	*uNR7q,9�ڬ��e3䘘�8)�����BR1���.I�\ڕC���r�ۘ4��)� (�xu����5���Hy3A�JU�z]�K�|6�l�r�e�� (�����`�s��,��s��C�1���#�Od���6��l����h���k�����3!d0����Q�Uh��j٦%l������	=��w1�qI3+-V��K��c	���,g]5&*f4c5�����֦6���ТD��k�? �� �x'�,��2�p�_*1����kf��g�6x�
��u���JO�`ԝυ� +Z2�g�oCӸZ����{`,L|k�����g�X0�Lz�[�('?���������8��k#�?���/ �Ğ��pȨ�d����$n�4��W�����W������������>mQI�;DOW>L<1� �V<�X��н�qQ�>?������H�m��q��?V��r��B�X�^��h��P:;�tv��捜����+�� �f�/�?���y��>�T����i�	s3�n���h�xq[����	O5H�̏�:�N�oF䱼�q��k���cqR��=�B��n/�Z2b���Z��0��^��N��QІPd������������7e���f���Y;헩U�ey�R��q�t{մ=���b�a�2Q��;̲��� �ݶeJ�Bw�ksT�ۯ�L��0pw�����5�g��]WɆd��߾��H��r�`��	�?l����L�����R:Ͳ�Zn���Fk�I��zo��s����"Lֽ4������ �Ÿ�łg,�T���G�4hf�\;a��¹�	���2eN�.I��!�Lm��������Ig�u�z�h��cJ���������jB�m���)�P6�h��BR�c��l�1S������۫���-���孅�hH%��)��Ǥts���N�;ތ��S���i��������r�[ �"Vbb�p��� S�&�F�i��T�Չ��c�3��5�"��؝�%u�1
��eD��.��u
��P�4س�b+��@��ϫ��O�0��EP�#���fY9�^{�� �hOF?p��Y�(�Ɨ_�V:ܓᰌ\�6�}K����W=�R����o�ߪ�zdH��A�"����/�16)������)��xc�'i�Im�c�W��s��>�^��y�;�-E�'�j�["��Z@x�����)$�\�p��!�Q��Qk>N�5��$����Ƞ�+���{s=����臉�M@OmB�ƾ��K�!~�_{�g�3Tx&*G����78S@�8i���>��Ih6�ŪCOl%�il�S������H��Z��{8��E������5��w4;$�2�k��؁毾H�W#��a� ���#�H�Uh ����N mԒ�Z�k�=��A~�ܴ����4���gKlT�z0�c����ʅ;�T��jDC���h A�6(��$���1��
�F`v� ��G �n���ێ�6�u{&~��e���S�����3�оlBRr�#��m���7i��To��DJ���ɐKn!�qɋ��5n����/X��|$�'��<����N�w�����۫�w��3�T�6��yj�+CM6+�"�"��á�,*��X��.lޟ~p�
��)i�|s��)D�x}l�)��ާ��y'�=���]1LH��A*��l�����kT��6���X�	>uH'71C�M]�4�����ك���0��V;�3�#�.�7�t���ff����{XG�˜KR�|�%}���c�Y�C�ˑ,��̚@�.W��1x�6����h�A�>�}�F��h�D/X��qA�1Y�M���ȇh\�D;|jOёj7��Quy.���^ä�>k<��V�ɸ~Ty��9'�L������Ug�yPL6U)[��g9�Z~�Ǧ�S��ʧӨLfq^�2�#µ滉��z�Qŭn���$���ЬȎ>9xC%UDS�_B�� l"��x�vz">�$�֟�FcU��иQk$NK@����E�l�q��;���K�wxN��t4*�xH����h#���_Y�Z���٨'�R
�L�5G���cՐܰк���>�����i.],�)?�^���&{���L��[�c��%���F�� E��c�-2ٮ������k�k'��v���G�5��@�E�L�hÇJ?�{ۤ㋬���:�/KpQ�I�$=DX]��+s�D�mYg��]��X#�iˌ��R2����<��