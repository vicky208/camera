��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:��r	��a������8:`��*ߋ'���k�J�t���3����Z�k) �D�}��5�����5j��N��u/M��y��	����-��t�푬0�k
+P���]�g �Ȓ��$��*](yu�.N-�p�M����B��EKv��Nvx�WU�@ƚ����#���]���ܿн�7JH)L���1"�ڏ�^zi��KmQvxY�#��0�cU�b� ��N�\avC���[����:-���:o�+!���>�Ғ+����O�u)�X���ې¢DeZqG90d�䖩O��)ܖV�Ӭ��oŤ�M�6��Ņ�1�v�V�;Z����柞]ϫ"�]�bQ椫�&N?��F��IF��ݡ\*�G���(Q�����r�Þ�����d��m�B���*W޼��B�[�K����r��Lh��O�;��.J�	:p����"/+ܕ�mMAc˚�B�� ns)H�U��������	��%a��]�?���|�h��.r���K��Qe��c��pf ��W),���/���9!K?SJJAb�k]Q^�.�����s�tU�ىB��.B����`�yx�Tb��O��g/$Z4�p/���ľ9v�2ځ���ֿZ� �u�a)<r�.E]�:�ae	����|L�VZ��
k������D��h$�bvX����A৓OQ��t>��v�F)D�r">��lxk�w�)�,������udͼE�=~�4D'��I�(�4�9]z�T�xƏ��M���t�<y	��Zm�*�{���U�)�e��ko#^B $u�y��BOmG7g��b���E�2�Z��]��#C��_����T64���f'�;
�(�d0���U�B���=Yz���o��/�Q=*��*��v��n���Of��h���V��V'��A� �uo��vm�D�d�_���k��늒4�1��[�����)r���8ˡQ�}x�W�c�/!�݉پ�9�w��{)l0jr�$\�;D8,^u����:or�NקK��TI�Z��]R�����5������֞#�;�̣�!��Xc���,(�=�Rj�ٳH�W��s�[7!��sV��[����P��@p},�d��F��@
M뙆Z���W�TvI��w��A���w��榔4��!|a��A�mA�P�.��lSK"f��)[���m��%�5;���{�J�+��,��.}���}�n��2/?�8��JE<}L�Z%/����rױ����T����s�O����X��,>��^V�w'q���m��24S^��d�������}cXj�Id��y(�ҤkW��t\�� ��9gfd�f�Ș
Z���T^�>�.y��U�3�����JL˱��aq�|����c��V5�!�����@��7CI����q��*��qy���Y�c��/Ʉť��)�٘�PrMyD�~�^����೦���ҿAAQ9��VAi�M���(p�Pl(c�ϙ��fz�z� Tz;
�5�4��q]2��Ө(k���6F��i�tdO�rh,��5-K��"����e-?���	�r�^�-���f�3��.��<�$�q����b1y�aGa
�V��6��>�F�Xא�~��^���0m�M@�a�]�o�~Ty�fH� d��&it,F�ͺ*�0�� �̈́n@2ge��L��E,AL��6{�b,E*�S�jG���c�_fo�E	� l	��\Q��i�>G���+��)ז���p�eY,�j�,$y�ma{� ���a$"sҷ*St�u�(�-���I�pE�vJ�yD4�3u��#ߥ�V&q�^�p5B񈑫�-ޜq�q�e<�Ĳ`A�*ju<�V����~�3\+?Ȳ�K�t�@�	�ϰ��̎�h2$��2:ZRS�S:�ߢg�(r�m�@A
��n�ߓmj'qU���È�fI�ꊸ��ȹ��=�Ϗ�Es�X�H��Tv#��c�ho>g'��|t�C߫�^���-������x��<���0�g��md���+I�B���:�f�*U�V��%��\�.��������W�ZV��
}iWQ���S���d� :ѱk�JVUh(z��ƎG��8NS�`VڝÏ55 ZY&�*�����U,�K����bs�"��;���*��
<T��ԗ�L�9�×y�oᴔj��)�$��l�s_s{�g�ܤ��l4S�֧x��A�\R�$����b��5x�9��e����s ��IA���Lr��D�'��7���F�t�3�� �v�A4wCɀ&��H0�`�ajm��}�`�d�tdM��u���|,���/���"+ۅ@/͹�kK�K�p�j�a��|�R;��|n�"p���%%ԗ���m������ �Vm SO�Zl�:�h�֬������?/�����Hl��o�*�9eOP���V�R|*,�ł� H�LJ�y���A\��R|g?�}������W��m�ԍqɩ�g&IH��OMMO�$���NJa0�y��/�pD�	w�r\�[2X&���O�����
9�>M���o�X)�D�	;���q�)�}ߠ�M5 �'�>�A�X>}���!�􅶠MS�_6S�=VY���Ș�۱�{%N�k��gdӴ�R��� *>�Pb�C��aX��mu��N߃��cz9�<�����1v��G.�p��M��ʔ��),(O�S!�N�������-�8nw;�:��?7�h�vc�|P��
�`BCJ�<P�)�b��F`��iT�F
W̵���tq#k"d����K��R?#��`��A'���B�a��9A՝4�ˮ�i�B�F��x�~LrRE���H�r����hF���>v	��r�0e�M;�'ϫ���������
���MT�	�<��<��f��Z�;�4�-2���$ˏ�D� �DT@&�T&�pb�N�/y��Iڭ�'����C�k�d(��?(3�@"���Ǻܠ���a�g�*��Ω/�X
� �a����N�[h��B]@�ی�c��4.y\cA�R���.���|V�����:|c�Z�4�����f�X��'�ޣS��C�Ӑek.�gph�%��W��Dg��|6�H6(x:� �~���H��z1�"~ajH�<��g��
R�6�r<�������[��Ѹ;��s�ݹ���=��5�ׂ��0`�2��a��ֆ�����#��i�LE�^�g�����I���֤�+��3g���PS�g��N�82%�v��5��PTV�(���N��^����2nS�7m�CCn�W��&=cO�6��o׏�UC�4E����@��8P���\O���S���f,{�w	o|	��ﳁz63m7�8�V�E`(��f�H�^d�P�nC,�Eo���'�D�#�h7�L5� ����a2�n�����J=Ql�����cٙx����4�R]�kbc�����U_�'��kɳ�Qx� �4�/��yi��[�4C_�P,�8��$8��
@��Z�&}bޱ�����,]�&R?���_ك�e�	�<�3�Ht��5z�\�����(.qA,�<#ʫX�1�)v�T���.\uF�7�J����]�Qo�B���<��p4^�/�ͽ8K���Q��,����P�{�s���J�p�li��LM��Z��ǹ
�]�O�Q]�"�/�
�n�ڴ�Cg��!�����5�]�x�x&�+-oU<#s<{F4b�A�0�B�U�l��w���<ٞ��0�!l�!�mځ>l�2�̈́�d���Hr���b���D�ˤ}���m�;M!��Z=�Pb��e4�" �~r��c��тPm�V�;V֨L��/�LHzoRa9x�w	������yÌ��f+�yB����]����R	6(�۳H]%���(�~�.��fAW�&Ǌ�w��!_6�lwo��c9�7�KIT��u�(�񽝲��|�U3�U$��MV��Ƃ6z����8�P�wݲ[ ��9]g	���"���P+�3�tR%B�{\����r��Bj薕�c�'�S� �r���]IR�l"�jLD&:��	���G۾�\�/C�O<�Z�����6`۴Api!��W�Qpz�Ո�`�� ��֍pPkG?�Ii-w>��Ne���QUUe%��wب��ލ!
��P�,��y��A��j��"APĚkU�L}�sҏ���(�9�J���א�Ob{X�&�����h���\C{�ID�� ����e�Q"�7~�.���E�/ww߅;�����c
g�(��[.HY�?��Ɵ|�T<�S�4�y� :u�N܃�,���rzw&����P��+:¸�ݐ��!�&N��4ԫ"Y��Z�Qq
� �h��H�g:,�^��"z5���_n"�P���7|��Y��R��]��s�Q��d���3�[�G^��Cۅ���0p��y��������ݡM��Z��;@G��{jr�=lD���s��>�v�}�� j��!��K_-�Y�]]�����	X�������*�Rb���(�i1f���Ӑ�����
*�~�]��MF>v�[�\��X��7��L�OҎ$�_�.��n^�M(3���[�Ǫ�{�v�k����J�>�e�@q_¤�&�ؐ�Rcv�;%9����;n����gs��$��{��^�ʇl��a`e�O����Zl��|,3��h�ɟqe����yX�Y�&�X�8��lR9�m�ŭ�~�0�	o�r�t�����c4:j%�>�Q�w�7�Ma��$~^]��p�ʃ�^R��'�8�b1�y~z�W<jV����)Hhr�Hg���Wc!l����;�.L"sP|��e��%�=(�+(�΍��_��9=Ml��g�~c�6�qXʞZ��M	7�J|����'�o�����z7UI����	H\Y����+3�ҵG"�j���h��fEk[dX{l�]so3jd�����[��t[�u���x8�	�َ���%�>�zJ�!K<��[ϚT�x�;������b�!�r��<�PG_מqr��#��R�B��W���_C����)Q4�L@®��@
��^c�5"WT�~�ܸ���G8]��;x��h��3B�x���k���W.\;Cs�F
bҩ�*1,a���SK��ˊ�eT���9�0ETLg- ��D���?�G���$9��eDA2��e#�&���l���@n��L��7��	6]g�R�b1�x���ۥ�W6�Ƣ`�o,�W�!�0����i���Ԍ�M4�؟;���/���)[��ף�k�
`��:&�f�j�tԿM�T���Y�� �۸�뜦�3�I�G��"����Y�/�/t����\�c��d$�u�4ylK���i�'�g�y����q�uWX�CI��O))L��"y/�=ﮯ��11��K���a�pmx	`o췭�p���&��4t/9V�*;0�2�זi'g1N�'�����zd_ ����w�!�U���|�~n�F���\\_�g�vD�=Sn�� �kD�-�"N*w1!'��x����kH �B�uATM�V9����pӔ~��!�a>2�)��w2��%�' ~㩁�3�A�e����l�"��~��@�<%��_]J��iE޿�0�`Sib�"������-J�o_�0#�#2S}i�ȥ��K�e�5}V�B�R��+1���!
ʋf>��x嚔��W4�@�@
؁O(���\sS���[�1� �5��V�iP�j"�(}O��B�+̟�hF�h�8�syo"�G"�[�R�<�F���	���ٕY"w^!,�ρ�O��ᣴ���zϻ��ik�=���H��Alfn�K&��Ɍp��\.%]:5��
�k~@�l���	��c�6�2є�9���������E��Ǡ#du��ur*��1���� �:.p%8Wr%6rToLK)_� tdY効u� ��F��˾�6�?�C���лS��M��/jva����8Q�G#�wɒ#�$��:���W�L͸�����%�,�pA�1��7��"iR׿P�6��o�X��k���u��F�73'>���P�V�O@�Q�L��(W4����&���h�e����� ���ګ.��+�~\%����?�d�P�� ܗ��X�|zH��+��+�[�)p��!)��HsVT��<���Ꝅ6F����lq�:���^Y�WIr���c���Ն�1D�z1�6�������H�s���!D�pVXx���|-�i����`�r|2��%�<]��%��ڥ��/�4f2��������)R�I��FkJ!��u���(.��Q�ӂcV�)H��0U����NE��B$��y�\`*��Oغ��1?k�8GXh���@�n�S ȁ��ŨD[�y.��������QÊ�8�K��ݵN��ms�¾���㖾���O���N�mG %\��8�@J���rp�8k�x��&�2�z�݇{1��g���<F�j�ډ#�,�$�
v����*8SFg_��3���y�ݶ�L�`��߷���H�{&:0��tm<Q0�T*��ss���O��8�=í�(����W�x%��>�BN�����9��=5|�qQӣpi��@��z�;�h+�sB֪o~�#���W
�dt"��0�y昢(�4���6w�4�����֝dC���0�t"�k���.�|В�Άh-���l���БA�BXk��pH�`��A�X{�^�VX�F��y{�{��D����R���\�v0�G6`��	t5uEF��$_��
@��z�!��>�`���%���MSr_���`���s�������*x�k�/.���q��R�FK��w˕4!���"��x7v��	m�y�9#�
aJ���������yO�:HCD	Ú�@�AM�	��wGJ2ܟ�Y�<��H�"[&7W���}0��F���`�<-���16!�4����z;6r�J�ϑ�8��%��*�p΀��,c�`.���~�7��lo!�2nϓCF��j��V�$�e�tY'O�p.	_�8s	7�DKi����񪃪Ҳ��?L�-�7��n7� �WN��X����<���cu�dȂΡ4iS����R�'�ٟ`8��5��8��O�>��m�^��"`FJ0�h-�e$�	e(��́Ղ�����N�9j#�	�������z�J�o8��U�H�0�@rKG�}N��49q/\x���"̊}������7
�z+�X��]��ZR����3�%��U�4�U�����6��'z��=�Քg+#��i���s7_Obeч����?�IAW�}�
�dJ=�N�Lh���P�JlpO���"b[;!:�ޡ�?�������E���4җ�v߻�H�\d��n;�p(��>�P�h��lݙ�\j4q�T���j%19*L����C8ps`�ѝ�5њ�)�rTAZ���+���'�b�]z(�&�,o/}��6�(�^cqP=}kc�s��,�[t�x�c�`kvf1�dJl�����Ɠ�]���uGI6P���?����F�A|^pg��,ҧ���ҁ�ҹ2N�C]��������M�E� A'��AeP��������`W�J\U�Ɂ%�����������9)�sh�@�v!��6����/E���u=]�[�%�9�6����޳5[�
1�!�����D�@�t��Bd��C�� �Z�()�雛zmO�aI�F`�v��@U���$��AsɣA%�h`R�f�5{���SÄ���P�J��]�{H�e�+��P��μ�E��q�(7��_a!�����5|�W����o������'��t���w�%=_��NV��6 �
&��SU�8���a�$�X5G�(��_��S�b�����AI���J�Öp�᫣+���KM�:E7���"��S׫�L!�
Rq��`�E&Z��.�.h@�����H?ڹM[k1��1�ŏ�8��7�����_����i���LH����Z����?����]�?���%��͐�bBv����wo�'���b��V/����:�s��̶�;3�]�րĺ�����I4G����Jd2��s 
��nF��RZ��~��p��h��{*m�T��k�x�+���݃;gp�F����/%<�3"L�=������g`8c�JԻ~�ՙs��t&u�$�5�,[O�݁�C��@Nѫ�1�M��V��j�U��߹rw��=�{��W�
g�^�g`�.'gp����c�)���.^L���}�CPt�@b�2ji���t���b�Ue�&����S}�PSb�!�GMQ��0B��a�� �A ���q�a�&h���٠�N<w����B�z#Sj�{�7���d~�c�������$���3����E�\�j�+�R��XAO��:� m���s�9r0�f�D��Y͸��K�E�)�z�IM��>�?
� ��F������QA�U",�����P&<�_BH�hq^�N½��(O�a��V�l����V��tv��#Z���!}�w�V�۝�R�s���dڿǡl�?>��%�,�Ÿ��	n�\��9AI��֚���n��i�b�1◞,@y�6��m����F�4�Z֧��Jz�2y�)��^M���Fd����&��w�7SY�3=��G��
-p#��+�$�gn�b�)����}~���߇d�I�KT�`w:Ǖ�f��bU���Q�)��,�fN̉Xׁ�Z�T4{XQtyf�gZ橭�Ž�c���{���g2����C%�;�؇�S]����!1����R�WgS��.���B�c�ګ�I:B�B��.�G�rf_��,�<���0��m�N�Vꑺc~�DH���{h;��sVu�N�C�|������QG�Cj {"}�w�|��(��S��S��0`|z[ԯp��/-y�v�4�4jh�̐�9K)�,-��MRc�<�?�N���r��(�����MG�AngA۱�
������-Ю��8��?C�aU�;�X���h���GG=��@�-ڢtSh���j�I�k�:a�f6�d��Beר0A
���lI!�B>�������ΐ��d�lm]�� �h�޲�OQ��l@:��t~�TBUK�@��'S*0����j1�.�IG]��+���܇��C����Q덎 ���Č�j���Dov����3�h�/'����ూ���,c����r&���2��Oƙ�8�)�A�s���S[�u}`-���<!+1f��mi5.�q�}�xR�P|a�
��Ӧ3w�DL����b_l"w"��p�����!5{�6�[j��Q�+;"\�{Ö�"!��:μͺ[�~��$/�ݣak
7����ڡc�(��h�q<���Z�{�OpR�+|n�R���h�mx
�9i����2��� ���)�o���㱒m���Pz��H����S��MbU8F� ��(0����1���hMH!Мp��*���t�Ь(�R|Vg��X��M�9����Ʃ�k����¤Z��(�, �_�����缗��FD��)�j
a%�4�͌{� ��O�����	��	���%���uτ�b�g�kR����h�J�ٍ
��@�)�E!�Z�H�Ϥ�k�� ����nx8W̓`��S��81�uC!jm��������Xt�{�)�sh�3��ж �x����v��e��8��tT�%O�y�S�zE�r֚��u��$p^��W{��_��[����ޣ����)f���<j�^V3�Jyi0-�a�KŃ�뗔i��E�K�����Y3�~?��]~/4�ژ�>�t����}+�� оk��}��0�@3UK�R`�X∤��1<�ܿ��=a��aX�f�f�%F����� �hj_�A�g��P��������b��e�~��~����HY�R,�b-u��:W�+���UQl���P����"�(�8�PȽj¯>�!�"�E�@��S��Dʕ�21d5�v!��a��������$h"���������i'�4?�5��*���~ԇ�"��1[����I�Q�������"�,E�P�/�1C�EZ�	���[c�����{��cǀV�>+vX��W��q6����=�2�9Wz�/���D-*�ۍBqW3^������Hv8H�E��gި8�܃ D1:ґQ0'�n#�NL*�����»���Y��J���5��|�'�v�E��ͯ:�d쁛�`=��T�׆�&����y��>
�Bԙ�H�oh�%A��3T��l�n���gO],gR�Y1؄���%����Y�$��T4��˻{}M�6�_s؜#��nRG����=x�L�D�7.ǘ�9���^���6�-@�������Z���/�ņbɷ�9t��Ƞ����:����҇<m�g�M�~���c�u.^�����{���P�k.��1��߭[����BJ�ւ��L��!�6�&�@�x�O�4�	V�A\����ZB�_�k�&�=f%A����Q��U_9�z���1,�T��uͽWE�g��D`�y�7T"���ܐbV%6:����Ż�� bu��	�1M���~ c�Q���N!�k�l��B�̈�up�Z��4'	���ep��;��Ŵ6z��s�Iu��>0�Rq�g�X��	-�I��,�� �|���i�P� <N�ҟ�c��(l�s����zq�n����-n_�Z��@5F2�x��z^�f}�
�[mX�f$��Rpe?��e��F �K�..Pgh�����9J�9!��)�jΩN| I�����>}�#W�`�*Cf�-�U������K����&G�\́�mdX�X�YGMI����\�X����� 0������F��e\#�;*��4��g�o{_E���2�Љ���7�F��bXV��-m�@#�!
��D1��Lg� _۶E�4�+w���KqSu�.x��\�]U��E��<W�)�x��8�2�NlC]D����Iq�_p��Ws,!b��%g����v:�|��f)�1�z���n��@�X�#Rg�V�8:��n�tX�Z���Ir��1��m�	�S����o�ʓ�{vr�LaX
����sq��� e�)*�NG���A��@!����i�ͷ�~�gV7B�m��R�M;/;�']�=&=���)T��hj��'��u��3��#�5�J��F���u�<+,&m�P���T�[$5+�R�8q7�\Ԟ5~'n$�pY��{ -%��}�A*y�����H�L�_�� �IC!�Ct���ߡ�X ������IF�v���l�m4o�g�X����xVN��iL"��	��߄=QeL�I~��O����#�����2z��Ȥ��#�d�_���3��j�;�������YpfZ�%����s$ �O�<Y�ž��P6�]5S���#���r���ۼ:���y'�ݒ�Wd.4��aH͔�v�Z��$�8���z�B�㺜��ޗ0�~T�:�[��xa������ӀCCM.�^��3@<n��R��!�����O(Q<2�"�@��BІ`�R������:�IR's���t��U�t.s�B)����������p�df�qT�h�O+g�a)&;����^R�:\%v勇���P�GGx+�������5mtHt͉��Tk��F�ľa�#�;�ڐG8�֭D�
�)��S5�5A�ʶMo�a���+�����r�`�O�� 敲-�t���Z�A	xI@>�,������P�W��nPpz�9����?�2��}{�GX����u/��t`3�&p&���n���JF7,i��x�V��S�1�b/[�����> �����Lԋ��٘�����< ���#0)���>ISz�X7��iT���l1�f��=~�X'�[8�h�����7p����d��;<�i%��l7�J:��d�m,mř �ntN�T��;|yY��	��N<ԹC'4�?f����H�O%����Y(�HC�qj���i%/x����Fr�ܸK w��+!��l�I��2�Љ�3���͉�#M��T��&C�"�o�U�F��!����F�2��/#�[-�xϛCC�]��W��o� �%��5�]@�q�Cٶw
��G�5��R��>L8�N$�l��tb�d$Arx�&�r�+�3�>�)���pO��t�N���Y(��#T:��m���}�NA��uOT=0���gk�J�W��f ��a-�sC���^)�E��x��H��놪J� ]��;9�y���E[p!��P^ռD'zh &��Z�S.�A�P�Gr��g�u"��h���{6�J@����_��l�C�@�l`���"BJGU*�|1���4\.XH3[m14s�8��_�+w-���=nP���ɏP���?�YK�U͏����M��|�:p�(��nn�;{ǆ;�(�i��.2���6�DUky��V���YD�����u	�9'7�b�1�_�䃹��3���n��͎��[Z�=n��U�忨��Dl�	�y8jwA.��A&e�2	<��|�A�eb�욌����R����)�I��]��/}H��NBCs���3ǰ;'�Ч�y�<1����={�GV	3�dwKO�����V#�]�H� ����q!x*K(�"~{i��l�DD������X���j�RD����Pr:Ah�(_��y�Q�sC�Mu���<�i��+�8���&���5eO�q�tWJ�J�Ӛ9��څ��<�T=�����ǂ0Uv.��g�mC�$8�:Vē�u���١��b<�A�IB⓱���Ba��\5��xK����z}ȶY+��0S�Uɺ��N��~F��82#��7I�Xݲ҂�+�M�*m����3�r��.7F~��`����c:��p����r�-�ևy��6��fJs���3�ޠ-8q�Ⱦ���F0�e�ٖN�/�#  Q�%��)
����z����]i�-��+ ��thC��8⛬��d໙7��K��~��#$9�9r�a������ܓ�li�"������G^���M)��*Wڣ�Pc�%�02U�CXS�do��/"I�.f�'���ʋ�Yu�k`j/c�����M80�����XՍ�e�7��y�\���hK�Yw��H�V3�������f�'�>I�X��hG܍Ux';�'�0�y��x�RDeR�[���X�7PN�\�#C��"jY�P�]�d�# {�3+A�6H��v>cpw���Z��`	��-t�e�#;��ha�K(-,�J�6�Z���8QmHҿ �C6�@�m���s�:�`�����lG:�@57U�*�����+�yȏ��<�Ā�����UQ\�,Br!��ف�$=Os��K�ȶ{���BfH��+o���>�+��&��$��ێ�J֔T&є���N�H�Tr��iΎ��)*����_�g=��4us�7s�)���l�jF�X ��)�Ic�n�}�|�E��.�Q9����`���pX�
��ܔ��줪X�%��٪t����ak���z�%T�j^�̶�Z�2(�4��� xs�t����:$�Q���!���D�t	!�I�1l�W����,�Qn?��R�5�Kn%�����!B~K�Y������Mc�(m�80�23����,U9<]&|�5z���`�Żn��;�������Ɱ�>�v�am�$M�0�@���K,=9F6�ʗ����	��.T{U�P	��mfY��,��d\��?��B���al����R����n�<,^
j�(U��*�7�y�A�ϙ7�a����7��r�H�@k7A��7�����2�,ܨ%�����W]�D˄�\���X4��2\Pn��T��8�<$Sq�t���@�E�h֮7B��8���ytĦg�h�J�3iQ,�*J��M� �Z��-�~���U~����"zD��m��Ҵ��8�jV�Za�����A���dc�C��2I{+m�l��׀v!�)0�$WP	&�a/ӱK"K�=`�f��M���M��>*�ŕ;�6c+���Ch�v�=W�2���i��˨w�DU�O�|��<����e`L"t�8*Ϣ��U����)�()í绖UcT���}�j`
[S��m�x���B��Wkä�.��eVfl�������1S=Uh�
EȞƭM�\�,+y �	�Zّ��j��6����N���RN�����Ecκ�2S/�䳟�I���N2�Y�&G�#<�|2�%�T��;�"E�����N4**(��-)\���R�|�X7�0��`��aL���	�{�V
2HwNnFmC&�[���@�<3|�Q�=.�@��&�څE�BsȊ�l(q_���:��o֘S�1�H���4�?ו��-����l��ڬ�]:�!E�o)�fc��12��%ܶ�nN{m�o��%�+*|R�gr�mµA7?޹HԪ�@�Y���q�(��vz뻙�t�OZ@Rj��ݦ2I���CJ)�lZV'�s�'��sة��	��xT:�0��si[�=̏���_77]Cz�l�h����0��@;%ce�:$y�
"詁�n� +w!�NVn�MEX������w�a.פ�B�YM?��*���s �w�8��EPg��&LS�z�� ?�A����*��l�4m�^, 7.<N�~S9o2��&��
|C�j>:�1�#����!��!�Ft|�EI�1����'��#ʸ������������߉3�A>��Cf�Pov�!Ԗ�<S�<�$RRp����s�+D�R?�2���AW�$�*o\W��X�Oh�z#�	%��4����Y�pQ��G��}�q�W?���La�Q�ʷ�4�X16�@�d��L:��û�\.A�5ݤW��b�c�O��l��s� ��$ X�SO�Ao��~�:�GTq����RT�'�����bAO�u�Bqթ��8~x�0�n�	�g�����d�z�Л3Z�m{�j���n^� }���cl�мs�����82���`�i�u��(>l�çh���;D^7ӧ�.}&��G�z~a�*��
h�%���|���XUTm��g���2.�f�ȶU��H&���+���N�<�8L: 0T���B�f\EOZW���B=�O��LP��2���ij䆪�@0>�d�����	2s2��=;"\I`�`G�0�.l#RQ
\ R+N#r|���!5�����b�d��!L�67w�N�����g�[�<�R�I�.��Ϲv��1������9����
ֺDr���^�����_݉^� 3Y�s(�5��<���kP�V<0�&��9�g����ܫ(���u'�Ո��%PMl�R�X�d�nm�rEZ=�+�i�N?����㊫A7�,�O;�

�����2[�N|�+����!��w��.�~�l�P8=L����7�L��Vh��L.>c!OUO��VDٮ�
5��LFߟS��f�b���{��3��yiOj���$�CXM�����
�ʥ^�)A�`�av�U�(ϝ�*���W�{K�ǰm�&�#%B�	+�](s�#4}���P�d�p>��|���Q��^�יo#ȿ̓�2C ��Ee��vZ��VoI��an���aR�'W^ =�]y���&� L�RF�Y�?�#�����xm��4�&��(�+�;�����Р�وJ��;ʥ�1$�[�S�0]�ÝS�Ύ�rΓV���Sm���j1`d��1��2XK����>?�x����� <��r΁��J>�;s�Z��O��Er��ά�5)/� 7���Υj��������xڭ����.����	�ڒ������a�L��I����	t?��M&�����!�O,~�y�Q��BP���I���t4����՞�P�c�*��$�j�Z�/(�e�Eg'��I#<"��V���wZ9�坻e���-�`C�D��?�3�I0������O_k4�e�H��	�7��-obf��܂a��=O ��|��N���.k(����W&����j���}�����@�j���YA�()0�A�+;@ҭ�/�g�	��Ƕ��u
�bmn0Q���v��O��u��p� m^�܍����*ȯ.�����?�?�ڛ\�	����ջ�d�j���n�[*��xta�M=��Y��*�XϺRJQD��P�u���R�����ӵ��qOY�$#�2RJ^	d�ѥ�:�ȷ��LOW_��b��v�S�I�-(��a$��c���Ij��5���,H&��1SO~�Ή~X{�氃����%<�����g	֊�J���τ���ͣG��?�,�xRz��{Ȭ2�3ӻ&�"�,gS���|�6�W��k�U���R	�@ˑ{v~w����8���ô)��$��E�y���z���T��[�?��Բs}�!~��@��~�9,�,H���qװ��ۀq�y��:�h݁�;�IX$A?�NKˑ�;0H	e�]�<&�B�����FG���M��rykN���ˮ�&�|�]_փ��b�&I��s�C�$�2Y��1JA
�uӴ�G�~�q��|��ą����(A�NL���K�>k�M���?<)�a�kCc���Mt��O6? ,�K4;ZL��AVZ��x��[��M�2c A3���Q��k߰���U�t�[7Ɍ���Phx@��K�\�!MT�h�l��t�k`�����Em�%��776)�O��ge��£��KMo��?k��K���!���ȱ���?Q����OG��
�����&F������Gj,�0�$�O�ү1�\ژ0*���@1�1�k��;�sl��,WW�p�ׅ�e�G�?�HL��dy+n�������y��Ȥ�S�� <�@`FK���+�1?ȎZDG��l�����r���<�T�@S�������~�%��g�N��, [�|L+P�g��r���d���������$���w��1M"P{ޟX�-h<��t��S��,��<"�U�8�RE�� ����[�7�تb�d�Vxb1��`XM���R)k��c���,��hr���Z���	7�����&�0]�2乕M9D��Q�;$	�(Tf�1k���5E���uh\#<��?�-��H4�{{R�E9�`~��i9x8�� ����ڊ������a���VMZj���,
@ ǝ��/X�=9�����/|�o]�m�Y���l3Mh�ZJ����5�'��.�lE���x"R�����w6�U�p���ęޜ1� ̅�Ҧ�X%�����ߑw{��S��fuً �Nu�s���ի�vA���;����w^��C�3��/��x���K�	\�#(%@_'��*rQL����&{�	�nu+���.�����������
 g�Ѡs$�=�+��-C�/:�� �z�<cաO��O����g���mcJ(�AY7��B�m�8�����3�
2|����$�o_ ��A�I6��P��<���IpX�FE孋� q�2�P}0f��j5�IrǴ��L�|��_����X��Y~z�<�>H�k	}��(�b�C�.�\�"��;�,׳K̮�#Z�x�4{��=C�O��{_���UHW�=�:*�R�����)�"�--aR��Y��aJ6�BD���/{�w�CQpO2d$�J����(��k��Jsy֗�0���!�!2��t��a���S�s=����l�O?�J`��·�(s!{�ΐ���򀿳�6��|��Y�(6.�H��ue�~�.�ɫ*�I�t)rᢩ�ٶ��Q�j%��.N�NI�_��^�J�QmK�)����1����]~�M=8	���Ax�;����f�2�齲j�� ����u��3ʖ
7v/��P{�1���b\�\OW�C|�׌>4���ϵ�������R��Ի�v��v��&#��K/8ҳ5����n��S��[�S[ayR�z��JyD�ZCf?��������Ue��8�`9tw�R�����q.�"�9,a/�yu�<v�}Ѳ�k�ˎ�:մ%`��`"��{���`����^p��8_�M���A2������Ê��)2Y/��MY�;g��Sܥ>�w��K?�	ykOD#�[l�W�?! �a�M�9wM�=v葬��`k�+�wP�feR�kZ;��ҟ�ʁ�t�h1:cg�0�����Z��
6R�+iV4���s�MJa�\JŭDb��cA܇��\(V�d#A�M�)�����:yqƨ�].=�C��M�]����l���ȹȂ�b���L�b<X�/�t=��sB�qC��T�|��}8�����,�D?>�JE>qd�\�����|�"��	 ���`v'ɥ�z�ԁT�s�Ɖ��7Ȟz��ty}��I�g��`�[�f?󽌛ӟ5NL���������%X吪:n��`y�5Ę��RLY�mY/U�݃�՚ �n���$��;�{�� �O����$�j֬�x�i�.��? ��؄���>�5����d�#}Щ�Y����p��x�`�i~�P���ڗ�ז���!�;���C��bF�%���*[�o}��kaU�ފ���Qf�bz�	��;�}��\�|ܰ3�J��9[+yJf��֨��]T��L`8�a�8J�E�אq�)#�"��{v�w٧�'�Jx+�B��.Q��<�X2�'xr�!9�N��ӊ��#j��Bqn���N������s�a|���5�?�(?����C�U%J��a���W�*Q�`u���nlv�'�����!;N�
�%%���N��sbs��S�N�������� �$!��U��4�2�_���/z�Q6�_g������q^�C�}Ĝb�Y��diJ�1b�T`� zm8Ȇ˦l�AbZ2zW]�+�W����)���aw�|���T~�D?��-���V��0�R���F6C�rzn\#��"iL.?V��$��=}�E���'�K,�_]��8�kI�^jS���yð���d����v�݌&��Y'R#@�l��R��
2,������n��(z�J�]ip�	'n� ���_����~1�#�
�_�P���u��[�r����8f�s^Y��C�g�䦴)�����(W�6�F�B�"�V+#	��Bo�����DIwj��S9P�z,ۙ�9�#�-������b>�l�%��׋ew�@fjߺD�Ï�/�r������8W��o3�os��	�y�B�����T�S��>=�����/�̘�L �&�&�x��������[u`JOW���yO��du���,�s��Z|~;�l����	�o������ZX�Vx��q�W3\�v����m�t�E��=�U����*R�C���R}D�9���Z�����%�֨�*:�r���š4n�[�lO�<Yą�"��b�3�-�ĢS�������N�!B�V" ���)C���3(�*��N�����/�Cs�Z�ѷ&� z(�	��,y�2]��:Z�z�U7EE�X��AfT���]����5���I8R��X����rܦc:���A��˴�MN�:a��|>� g�찏Bw}��G�Pzo7��:;�`��Ք�.7vn��M�_x�"�;�@)���56&�+�����-ƒ������"<�X�j7�2�Ӎ\X�L��ʝT�����л�S+�M�Rx�U��`Z>l`}3�[�#���cz����(YU���FF�w_��u|���3�?wx�꤈$ML"���&H%K��7���{{!�7/����X�$ۻ\QƲ���}�����T�Ml���_���Ē-j㈰[[^s�F�0$=�.�RDC���v���"%P��7�T�ʋ|��ȅ�{�X��EU�"M�)<�&�b�@���樕B��1��y���5�#��R���'B� �8#��?���w5��k��r�3 �,|!��q�ޝB�!<�����?d(�$�"@؍`�nav�]ŝ��*��4�P����F��ꎭ\�'�U���R͕���p7��z���;Q�W�9-�g �;=�̈́��y���Ŏ-<�)wrّ���dㆦ�3>Q��"��My?X[ �"=�lw�т~��>���6��(�eK[P�B��p�Tj8�h���M�{Шh9:!?�)N"�b��3P�p���H���NL� ��
^?%�����[�W.ߑ�?K[� �Ҙ� ��60���|����_� ����bh
���j�&��dH���n�)a<=�mn�����g����{�85�b��/>�+Z=��|ж1ܣ���Y��V ��%9F�\K�ޗ��yK�hUB�f�!`�9ZA�e8%�\���a����Ҽ5,�Bnʬ��� y��� fU�N.K:)��po�엊<_��&����P�pL"1o0��<=��(��k��� ����b��-�j�>���C����@�w�}�#��˘�1+��/�Ks=��.�=*�q���*z\�+?�X��A�������d��*�Y_Y^YkjU/�8=�w'g�%2� �ػ8��Sٛ��T�(]u�O�V����wL;m�=cς@"$@8L.S
^�]\�
��h��gg|�I���;���,�@��"�ǩ/�W���m�8�-tJXTB(Pۅ�_`���2�L���q���p��C��>�/6J��
����1y�$%���о6�_.�������I1�3[?%U�1׾�cf3�2�Gg(\�v�@L��w�`��#`���^����>��a�l���p�v��Ю�O9���R��g<��@\�A��¤ehw�%����52u���=l���u�������nGש�Jk  Qx�0fN~e�9�km@�0��-�;\fmj�}<%�{֏�pAe�Q��u��J7�p)x��6�4Q��!�A��$H��uw�s���N]��ڝ�^��<Ow���0�T�ṽۊ���C˂�efN��˙P�JEm̒��K��8�D=�x�_[L^���Жc�e��vx�.x���#/���r�l��2hL��e��� ��T�?-E��H~����Ӓ'�C�U8 /8h�V�d>��w�0��6Z�3,��I6��~!�%C�.��~SгXrAb���	�j�<!] }h��O�pU��Cu�T�^_a���D�:X�����CWS�ā-[D�i��O��hSW���0��E{�����[�P�F�彇��%����̍	uа������ҽ����b�ޑ�CM�ߟJX� %(��{ǘ3�$�R8�R�O	E�;$�),�� ���)2KG�x{)��1.���f�
�|�61��~?�f�~C�b�ixJ�6p��.�����`��c���|�;�[꣖:DS7gQ�H&7��	xD���/��wy�c�S�S1k)~Y� ��i�	V���������Tz��Ú�r�w�뺆��P�$�-�6!��U�����dO��i�g3T��6�y�Cr�:����Z��p(�
�w���i'W<�����RH�Yׅ�OeY�d��A
.i�p"o0�����/ʁ�y" �ާ�91��:"��B=�_1m� ��`0�"/���>XG�'x+#���Vt��^�)Y�+:@� ��" ܡQ��E��D"��I���}�J
�B
���od*�eMg"�[�a���AJ©E+��؂�����{_p�*H�*.�<�1�<db�N�⚹�@�\���5߿����D���v�k�8(�P��h���o�]fَ�ϫ���F_�I�����E\mo	e���9�ύ��h��	^�:��z��h��ͼ_8�<��"D���4@᭴wR����I�k���������4�`�b�b�	H�'R���@N����
0J��Y�nYl�.K�����hs�<�� �v��$�*�E���l��qDE&f=���)L�/�(ۘ�M[�+Dk{P�T	�6�{
e�����Xϸ��	I=.]-���_��,@XY$ 4E��:�yNT3B��ܜW�:�rG�d��pi�L�''Z�R��$�b����4�ڕg�	=4&ӸCǉ��j5&���'܆3b3T�$�fvSB���W�z
 Y�c��(�s�����%�Mҗ�P8Oܶ�E�l�K��vP�Ԋ��_+���5Ux C�gOه���Ccn e��n���t%��˙��NqvMW��V��ZL�W�3�Jk�X�Z�Ӝ�5f��7_�
�ƈ�+�Î)�̠�É}����R����@ �3�7u
�Z��r�s���s����)	XTm(����b킻�-��T_�`��p青�$���_]�"'�,���[��0���؂��e�0keX�4�T}�N�Ps�|�8����-�EbB�0t�O�ci�|Y��8�$9�dn-U�e�p�X�S�z�_����^Q]r�I�CTбvA{~Ա{�^��5Z�A����I���]�8��S5���K�:�v��S�R�AM�0��0G�e�j�\�J`�*�ܔ*�O��Ĥ<�&W�.��4P����tR������dB�֭�b@űIDM�o��t[�aT�ف��'�ʈ$�H�}kSR,%����͑�w��T�hq�p�04��q���@r��&�$.�����;/�	��MX������->��<���BxfDT`-�>�u> g7�Y��{+䔊�m:����4�:!�KL��g<�N�� W�9��M$��F�Z�3n���'��~`!iy�qib��K:]��tI�+�h�[*�=�!L_�u@`��}6�Ŝ>��c�a��/c�3��$��.
�	��}T&u6��M�e��S�J�A�qj�	-�r�����+��(K��qf+�w�؄����S���9`�$/Y�Z�8���x���8o^�T�����r7CM6�7sܓsD���GH�d
��*Ov�QՕ7���G��G35T�qn}pې@����~w``�j��,V���.�X�=,��_#��Ꜿ�U�M�`��&��rf���`p&�Ima����0?��K���Bp<�¯��ܦаh$ԋ#����W� ���3m��I꘺��ZY����ΐmo� ���抹�`J��tΏAnч�m�%�� ������I��T�}R�h!vMt�!�G��l�:��/4��#���es4H���|��'8nv`����w���wW��XOF�)��Ù�{��a�o���x��%��)ϖ,5�"���n?�f��+$��w�NF�r��!�4�Q��R���{^�����>wpRQ�%?w�WQ�y�5"��gu��X�&h��']S�ƺnT��u�p��x�K�d?��H�{ne?�BV�"h�$9����%�Yk���p�	݆��p��Z���
�p��G��%�-�9�7[%�	l����8N��KԜ���Һ�DW�i��S!�r�aT�>�GKpn=}}H�3��/X,"�a�Ӥ�I!qS��,�(��F>	��f��ٟ�d8E�G>�-�x*��R9��Ed$PWt�:K��<n��zE	(*��9��s�)��Y=���:P1�u0�M�=�GZ�O�Y=ز�p˃�N̔
8�@�Ȯi$���Jx�Z9��e��m>��Y���� ��O��بmoA4�;q����Ek����������%�a3p׍S�=K�_<�![���Cg���ߙ2�qC7�9?���~i��������F�L�v��wkL�D����b�k��Eq�e��i��e=�&�X,���G`'I�� �`�9�����к��ӧ@D	��rp :=\�r{ɴ����T�������"k�I0N���w#����Ư\�����ӧ
�F,���vݠ�V"'�o����C���X:�C�a������a[Q�H�%E��H�|�@-�r�u�����ᱴ�pؚ����m_Ҁ�ˋ�UiT���AU{R���}(�?��6��CHD��R<�P�_#�6������3�;��뢹�{f��S75A��Ώ'���tz����3���Q�����i��'	1������u�^�E@A��)����
��r.-6�+�S]BU��?!C���f���}_]�E`���^�mG�O18cV<2��Ο��#A3,���6
>r^����dĘ!<�J��~�:}�-VEb����\�>���o��H�����X���ˈ�~с�{�PWe���b8�^V�\�~��D��(C-R� �ݤ[í���w��p��3L$����q��4a�Eu�����1��[��Y����pg�\���hV8�g��q�E1��\ׂ��S�,�.�_5! �&qt�R;wuӔu�5G��S����}d8�7p��8SM���\��~�/5���^!�LPe�!�(h}]8�?J'a�-:��P=�t p�պa�$��ry�8��M��,��ƈi=6�i��}��	���3���];G��%��a#��9��O�m�W��`^]|&��|�'�Q����w �$�u.�B�"�|6��6��ʤ���!� X�u��y�G1,wܜ��z�t:����R-R%	���2�Ƅ!Ä ��R�)Bz?��'�*�n8��Kk���r!��B����?���l>LH�b,^���G���'�G"(�ݬ�\Ch����V㍛�'�`���Owm97������rD<s����e�\��ڿ:��!Pq�B���(��R�2�q�Ck}�.r�i��g.']� ���<R���8C�k����\�
��}[�}���, Kr�,�3�Y:�q����f���0ī��'��|�a����!����kU�UL}�*�v.�X׹�uQv����1�Ԁ�YX-Ͱ�dVҵ�.�Do���r$S|,��Rt��ڼ���'�q��%c���f�R�fY�^�z��ꒃ����T��+k�<�-��c��rb��B��Y	�{g8y��t�^9.R��A_�s�(��{P\|�߄�=�+�>S�Ŏx�����
ϿkS���R��<���W�V��!45P�
%�(�:���?��S�ܟI�G�v���;�
�	�X͒���M+ ҭ�O��[P�9ا9�ԍ�[�y!�/�Wy]3c"x���y�CY�,y��Z�fW�R2�2^b�M=2�(]�E���V��PL죁�¨[D�(��r����ٜ�/��ý��$��\� ���������H6�\��g�t��PC�W��U$>@�}���ϸl K�T+��b�9F�gl9ɵ���P۟W@�f)ߑ�A������DC��ݶa������`������.]σ>`�q�G{A��ju+AsA�:��-�X�zՀn�F��o�ɻ?��H1�=<?i���㼐�N����ȏ���fs�(Y��cJ��q�ώT���ͮ��F�lQM|ֈ첪�2����7G{\RͰ�[@I�S�y��7�"��H
t~��cl��D-�®�c���qH� ��ynU������:�HՀt�|/�Y��>���fq���͕����~���._ȃAĿ`g�!U6�������I�Gu�̎,�8
�^��ot��ܛ��נz�����==yD7���9��S.���]�J{:�D�� 	��{ͩ�w��a  bIh�d*��f*3����ǉ��]����*�9�CY�T�|{��E:_D��:R͉7���W�!p_���|��#�6��o	"�3�I�\��ډD�P�4t\4-�?3�6\}�DvH�b�\m�sƿ@��f��#�_v��H��y��"� �j�krjZ1w��pR�����؉��+�*�6�2l�B��/��nDg�P�����|(��8�!cvi�!��)��_����^+;���18�5[[*�Y�`�[7	�Ȇ���H�̒s޲��U�=U��DzW+G�����`�>��9���>�ܡ �_��8e�#��kІ�ϟ��Ţ����|i2�1��uZ(J��sW1������=q;D��@�`|�Y���J�o�s��Fx��=��fp�!���9U|!�yS���ߔ��E�M��l=�D��jYϋ���hK�����:p�<"Mb�l�5p/����2����6<i���Ҕ�/
jK��z" l���x�z3�J�o�|:d!��1���p,"�[ˇ]e�3���<*d�Q؂D�_�0y)ޘo,���.y:E�R��T��D����w�]嗴*g@G2�!� �5�e��t��w�b�-���2����߰� �H�P�)����q���Z���q�J �7��%���-�N������o��*�㮉f�N:�i�{�����������_OSc���m}�a�	��+=�6�Os#'cNx�����B���� � �Ƈ��ʔ0)��|����E�[f����dg�U���HP+�|���N�&�󫷅;A|Ǽ,�Io̻�g��<�5n�<$L�'�׬��uژ����<��kh���:{C��S�����.wV�k���+Ihi>S�k
qc0U��ũу�L8b{e|R�i���f9R��m�>�^�p#-T^�&������u��/)
4������Њ�率P/�2"��!x���]�R]0x�ZL���Io��ڗ��zi|R�b�Y�4�[N)M˜\�b�-��L�i���2�^lY����b�W�{z��/(��,�5Q��j��G�
�kl}���=�tdf�2��Dy�,pNw0�xƂ�Ӌ���x'.�O��z�W�}��n6W�2����lޚ��uK�Li*�ˀ��~c5^Xoɚ�"R>��I�(�T�:#6Я*4�I�}7.K*ĸj��#Z�X.f��y`�%�"��^�JC.�ť�	��Z�\�r�)H~P�?��P�G�I�,�!&�I�ҡϑ�B�<2��ؤ\*rz�3�v�=l�E�$�*�?� "K�	�9Ù��lWj`!���<��5tX����D�!O�w�ꪪ�����]b<g�wO���?R+�����xL}Rg��-Y6��Sb���N���8��s޵"�ǐ���d�[C[��V5���א��K��l(�.C��OUl3���
��f�T,�����������#[4�۝e-8!܈[� �ׁl0�_�m2"E��V8���=��}솥�����Ǘ�#+�T�t]Y��R�I�`l�Ȃ#���@L���G;Ó�� ��#�C$�k3�B�r��G�����WJ�q��Rw�lC�d����"<Ĭ�7�z��Vl��q�y�IzT��U������*`�g-��h8�E9���O�Q	Kہ������?$��?��8�'"V/�C�� [R�b�<��.�?�Z�ѳ�%R�K�l�xy	��N�Д��}����2lC���6�"�K�!���O���k%��f:��8okFm��~�
_S�0y5N�6',�D�,�a���@��2��ă�%Ҥl�ɷ:�H�u�:ȴc���^-��O��B��Ň�JN��ǩ�>+& NSu-!��_�(0��7JC��́s5��<^��:�8�A4��&��e����l�{W����o��Ge��KzoЄ�Xd8Ed��s}�>�m��-]����m%ϔc����ĭz�:����
lN&O"�aL/����p`�>�J�Ӽ}�I�e\ �I�<�e �9Z����ē�;%�a�������� ���`����������2��9YPq-�-����3�� O�n������'�O�-��TC�����S�m���5���<�@2�۽�8+6�ؖ26y�8r��
�o�{%G0��,�^]<*�<5�_.�,l��UzXR\���}{T���7���n��U��R=7�9����B�+��%ƛ�O��r�~O8�#��HB����Z^��w(� k���=>/<���l��2K���jLi���C�[T킚w��.�\%��)��`/��65��=I�j��߾k���@lS����߬���TQ�F���yc�C�Z`8I�<64K���bDCM��Ҽ�*̷ƹ���#�4���rC��˂���.kOЁ糩�2iʁ5�_H��|��j��)����1i,�G[�A�'�pp���0�A�G$@�.W�,������.���hs��M�E&�X�f�� �(_�	�4\���	���S~�EX�I�Κ[�:?�A4�S�Y�� �_r������A�|�e���+o��u8/��=>d1�UX�������&.ȠS�z�wL�5݊��b�0�1,��g_��֎�[m�� 	P�06q������<w���p(�$���f�B��[�->��z��AjP���+.�aa�>�eŢ9�Z�ӏ���=>{^�����4��i��°����=��<�"&8�m�<�u��Ȅ��7�L>"���3�8p��*���K��aSP������#�e��'��l�,C��D�KÉȤ 񵭭�m�ߘ{�o�V���g�v;L
�cWJ���ƛ�=X��W��������L���u2�
�?��$Z�9��l�����8"�!�`XQ|�F!IRB��+K�1�(��Yt0����V�S�s$8�M����4��*����]Y���20�X7�ލ`�
J�� 7E
�0f�	^pCf�^�t��� �T���1jUD+*8�i��ڋ��#��k&����[��i���3��<�>�ki�@̀{��2��0F����N�``�� ���{���z>d3��e�"��%�8E �O���A)���5�H_n}�T2�1���V���:�����Õ�� 8����l�k�u�gT�uEP�=�gL\��G�H}�����R�z��=���\�[���Y7�.��-Z��Z��]v��W�j	S,��
o���;�@-�paEw���t�'8�FP&��Q�|w��>j�[O�`ua�S�Dka�Zv�*��9�h��aIOG�"�ѻ���_��.�%�T��:9�*����B�[i�Y���>��`�Ro[�Ri����{t&��+o�L���G�^����cE���-$,߬�6Y�y�¨nm����R���9yS��#̺��Խ���Sd΁ZN���5E��>>
�Aw����y鹧Lˀ�*���ԵX�V�	l�i���{3$obu<_�m(��'���E�գn���m�i��Z:�QJC^/Z�n���Bݭ	LN/����@j�2�N�F�(��$�'�fblVgV�`e=��N�����i��~wX"-x�������a����3I`e7Ɗm�Q���+���X����˸�/�ޯb���o,ܣ̗��s��E����{��;�����ف	ެ��j�E��Ua(n	΅\���S�
)��#�H�q�Aw�� ��\�����]�Ga�m"���ϕ��6Z� �u�$����Y�#��j�U� G�K`�����ȿI�Ǿ�V��鍊E�q�:@�N�E��~$oO�t_}#ߵ�^����w\tË�+�����a�J͠�1}
��^������2,T#����)��7�S��g����j���8�h߯�J�b#���_n+���V,޶�%:9�@�`D�Z���w�÷6$��&~�p�>'� 5T;߰��۱�C�ή�>^�Q��� ��ʙ��y�J��l���=^N�weg�꟩g�l�~����N��0��j�8s���q=:�#����v�|�Qh�隗F��zȄ.%Mw�I!�9�H.�kɿ������cXw=�U�D��}�F@�����DT�Č�z<ͬL��8�q�/��b��p���:F�W�.q���]a�U:z9�5�޼u-�~��o�"Vh���#���;E��Mψ/������ B ��ΌjA_���ΎԵX�+}P��Ml)�X$�a:��q�z6�|������-OE~yH��\�l/;!p�5����mB^�T��=`�x�PX��B`�r�:�2b�ު����"ܱ�\���R�dc���$�������ɸC��)��L�L!���9��WSJ`PR�A��_E4�ou8ɣ�DT|O��ݤ��6�n���R3V CSY	Ť��-7U�Ϩ<���ۇ��!�C��רlH�NQM:�v�/��5��EޏER�`^�P?�'�����ȡ�7��y�?
�?������q�GmY��O�2�c����6�pc�k�Ñ�����rS�*�����mac��;3�g���Iյ��:�3Ś��@��Z��ݷ?��g���A�r��v�Ua���Դ�d��G9u�)J��x�O�S���!�7I����)RP����������I*`����m�Tf0�����Tj�6�!���1A��G�=8�^ȐF !oӢԣ�R���YKP�Ǘr�4g/vZ9VIMm~��|ם�q�V�MT1���!_�%�X�N�;�S3IA'���&���w���^��]'�h-�'LOt�����t�b�7�[���?�u���=��Pz����,3LI&�wP20�{RMx�������b�R
���׎q�2�:"M|��� ��5h� cb��.��rٳ\�z�p�7�"݇6�v�4��h��J�>6<'r��FZAM$�S���3���N`�D�����h�[��A%'�l�܌e�Ʒ�8�a