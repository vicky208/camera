��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V�h?�xrMIp*/�p�x�_?�F������j��1�v�Y$nq�ˢb�=ᥦ&Fce؊<��������Ƽ:~�I1���$�k|X���TT������>�')�>��<�� i�XA(~�%�#�r�yw�
�]�GȺ���.#��K���C~����#{n��Uh��^@���b�"�2,�Hu�
u�x	��)��0|Dvo��fh��*�wr0(2n0��ֹ`�N����:�w�s�QG0��0I����`!��?�~���9Ӕ�6�ݕ�~ue5c&�Y%�o=s�Շ��d�ചl//��5~@��*V�6n��Y�"�f�8���mSb����ê��:鞲Ӡ����|��/�"Q�@K�f���.�Ǣ[��#}�6)�3�^���7�)���,��!�Ν�@�i�4-:�x���i��]W��\�t����-�@�a',�(ct#6�|z�j�0�偨uŴ8��U�8��Fr��l���Z�Xh��gI�l�s���C�p�T�>qPڰ8l>Y���2�a���A��K�O�9ɻ�ua�8c]~LՎ�qG�FLd�F��W�)��c��/�rIY7��-��B^�D~"D~����,3Y |�h��}-��I�_��T�_ҋ�{ �����5���Ӣ�K<4ÜP�U7�����!���x
��l\������اF�+����~C$�����| e"f���������W
}����z �Ҝ��������%�cxF_�u9��ހ��!r�}8
R+j��^
�z��0���g�5�wť�̍aq�e3�A��
�գ���[��B�CxΦ���5m0�9�hM��߇n��q>�`8�2���j��8�$��f�?���Q�Z֮�:y���c�4e�<����C%�vRG:B<���7���}���.iţI6�о�b��������s�3���6������&�zH�Y�9*����K�0�-��������=^�ot�t�� ~����d��G�ǖᐐ�7�{�\I�U@�AVF������k���?w�1n���ɻ[�.�M��+�_��VZz��<�Z|@�J��F[�"��*Y[޵Jy�P�����AYjJ)LN��/��;�Ã�k�/K��u!|�X]Q�
�^[
>Kp�nxm����i���s���@|E�ՠ>��X���{;:(���Qé��Y
be�?��u�n�ۻl]u��H�iL`�5p�V=�p&�l��>���Mֈ�mZaL9�_��T�m�|�o�(�JC�,���Q+S�>�z��X�ݡ�}���b��݄	����YZ��������܁M"��\G-}�}�MHh�,^_@��$+ۈ ��1®�8��P�C�6{�'x��E=��Ri!ض�IDQ|����!Q�ܖ���	X��@h�w��b!�a�QXV���rʒ�y�!Rv�0�������{��:f@�D�gk��5�j���].� �8l���.C����T6:9�1�WۦG������g-�K��HvACO�Yal���٦�}]�2$^'����VRY��(�l!�8��O!F����å�����:��tw�Xͦb6��/�J�o����)�MW��6�9�Q�U�GM�$�%�z�iz�����q ��13�k�Y0���T�5�)8��'?��6`?q�ٖyB�h�(nJw$+�Ձ�nM�]���8��+��BZ_�)k��bMUb�d|'��J�&��o���O�o��ɀ�$���z���tc�����\�no������FITބ>� $}6O{��`Atq���+�rh���3�Jx;�+` ��E笍I�D= �l,��'�H3���!n0WGd�i�_n�E�>c��(,��{����\�L7��Z9����/^y���%�l7�:�V�<ϐm�i�́�e���RcR�u����q�Dk�=�ZE�
~���M�c��r�|������XØ<�B���<ZW'yۥ9
���l� 4�0t!Snݯ�$ �,&-$f����\4�<�O�4������{�F��Qt��͕�e%Eae�dڝS,��h�S�엫	�9<7
%��|��E!����J��J�����L�U�������j<To1�7��`2���������9M��;9}P�����^�q�&��E�hsc�^x����g�Fd����1�/�b�D1ZsZ�l�`4�r�ʴd2,UY<��=j1�2��j���7�Cyy��E�)�-v;Iǵh�U����T߭eo;)8�_I8�>��QB����Js���6����J�oD{K8dѭ|M`�_����l��N��瑩�o5�9��>SX�\�vh�hb=�j[f�`#~�O��CzAC/��N.�]Y�c���5��[w�<�54^���!a��K��ugdI/I��>#�Ѵ�zX��&YiQ��3d�@=��l|A��E�{�9@�I\2��)#�#��Y�S8��l��t�e���D�Ԅ�- ���g>PQ9�$�_��8D��@�����> �L�W�E��;d��@�O��������*T�W�sf�b�f�K}K�Y� ��ܰ7����F(Wd&eTZB�V�(RS��7Q��p�\VQڭ��1�6�]��SH�u΃}D=�vр}��P�W�/�1�b�Q1��p�~瀊0	�؂TY�:�4y<� ����?�4����q[�Q���y��}#�n,e�.k� �4U�'��r�Q�����Z�v�	Q���0%VZ!VN��XT�ĥ�%b2�aU�������U��5�̎�������(��JD�#�[�A^��
���7����!RV�yЛ�o"�|���W�W�md�U�1Dk�Ҿ����tCX5h 4�`�PuK�Vbv0�Α�:�+�iq�\r�ڧ���i�.���K	OI�@�Cy��R�"
t�yf�|�	�3n�n���A���RwI�]�$��ߔq�����ލj(&��� �	�.+�Z0r��巒�OT������Z$�;�,�
�r�}ro�d��2��r9VA��b��?`�@b]Y�+�'�p���4%�l�E �Ϯ�8�`:�-�\ll�-�O��[�V	LyT������X��(G����"�@�\ٯl�G�5C3l�!]`�[�AC�_��Pt�V�_5/�6G�[Cl�0ꨠ�=�c�t�F��!H�����+a�!1|�b���U�RY����U�q��@�?T�q���Sjj�^�^�:Z���ȿ�N���3e�^�Ns)\��#1!��)�B���W�gr�o�λ�Q3%:�]&��*��S�JE�Ki�qZc�e�a���ν��A��u_��t���7г��7�n��f�4�''kt��p�Uw,uD��7��"�������ۡG+�)nsTH(&Ǥ��3�˪w/��<u���4u�e���w"��mZ��b�	8��RJC3�;j�����b�����t馟�c�.�r����c*�sE-�Ӻ��u�&Ϳ?�{���\[�5��v0s��#��t{)�>I�:�)�$U�FSb�^�f��*����?�N���ʄx�@�xY�Bʜ�i��h�/�r�k�_��?u��i�y	�bL�z� �#)j�V��<��.���ƗgL �
�pA�Ӄ�}.������*ިJ�R�j�"|���\����?��E���Q_��!���͜S�\��`��*�r��µl2��(|����DS�4��D-Zh���ӧt��>X�,��'�ی%�m������h)=�n�����q��a��5VOM��Sנ��|�C�Oע���̍&�q��z��N^J�x�
��܁a*ay��t̓��w�dWx_+�]$/c> I�b��\�r�l����Xf��x=�<ba�UR�%"����]��:\i'�q�E��<����ܬ}�c.!�����
U�Δ+@��v:}ê���Qw��X�b��$2I�~.�ߙ�d��	��n����6
�[ ��-���cE�n��˳DA[��pb�񱱊��00kx�k���]���_ ��M�'�g�^L�����PR��)���~7�̻B�pXjϽ���7+��^ ��R�jhl	���W��Dd����	c(���'��r��AGce2���O�A�xsB�+[F��d�K<7Lݷi6������<��A�&'��n�\�U@�墏����M,�m.2sˌl�:6�+Iz>��X�m�qR��z[�;$��E�h�����1n�a��ʫ�����!�MD�i�#$�8�~�Eڏ��2�S�V��#h��?��J ��M&�e>7͂�:��I�j�ɘ�9��F%��k����r�_�ъ�ʦ���TRŋ��LŽwH�E���U�&�Q��QӺ�2�,���)2m��gW�`���O��VPZ�m�6>�~s��:����E;����O�b�B��JSN�3L��錣$��2�\ˋ�:�7�X�S�L��{�$���'��Ć���[�Y`������*�a�����Q�w��
<z�r��r/�ݾl	wI���^���wcj8���(J+�7RfudLQ�f�5~��9o������,���pU6+6Y��?C�͟O�	�����w�{�,R��B�_Ϲ��2-\%��j:Y@WN#k�����_���$��'�!t�A���C9� �*��K]o�6���ϑQ���� :_�ٻ��#�E�6x���Z���7c}:����a�7�����o N����k�c/��L%��>|�aϼ�=$�����0�)��a�_ >��~�د�*��#�
�PXOm���e���_D�-ޜ�g�0q��U$���-b�,����$�9����.�V�l=�z�ޜ�Õ\ �X$�i��9j���l��5�N�q$�^��*���lm�[�ƒ���kN�f;1�6r�Es���stQ6f(E/nl�٥sGp �?��f"y��Z/�I�f1�	�mƎL�.���ά���0�$ڳ�F��0JW�G����]�y �;^�A
�=�Bý�-ح�w2[$O����#=D���"/Br���$'�Φ3a"�9� �h�ɯyǠ��5d���_[`�8ѡKid��4�������o+�,�Q�:�|Wl�b<��:5��2��|�������+����W>K[A�֤���P=k̚�յ��H=5*�?|5}.�6tY���i5}B�٪�Rڑ���n�rOS�ԛ�5X����eܸ�2N���%���DW�AY�pa��<� BS�/u�k��a� �N��^8�ܺ�P蝳cc��+P�E
�g5>���k�a��U`��0�/G5gP�"Ʊ���FR\$8�� '@��?�f�����8x=�z�]�'6��nT�:�A��3t�~u�Q�&XWR�XtX�M�<�U�XA��bŘ��lz_D�.��3��a3L���K�\S��Qn(��P±��v�R�W]��n���m&���
�Of5&?r�3նh��j�NU�@�8�H��pUo��[.x�$YY�Q`��8��\���n�"�S=QM���d��r����o]c6�$�^L�F�����p�4'�9EA��YTD_�],��#E���2�2۪��m���߫�c�0~4��ܮ�A\��/=V,�b�t~��C�u� �o6R��9 �J&�μ�'L����C�Pt��" �Y��V����L]B��Rۈc��<�Ӻ�wI݃��C�����O�5yt�?�:�tO��6���ڕ��߇xw�䥙�%�bb�(zJ��YP*kmL�q��Ђ3�:$��m�恑�!�Vv&YNk �:��1�F����e��.X�X,�ݳ�����VJN����Z��0�E� AmѾ�25��l�ϳ�j�,�T�X�S�Ë5gH�Pe���[��ɗ?!��ŋ�c�M����^���~��E��1İȉh�2��ʗ���H�p�Aw��VR��uU��`
�hl&?]�J��*�0Hp
�b4%�"�~9$R�w�<�x�ӝ4�FM�a�D�;��������+B��rX#� ��?C�Ѯ���'����=wՂ\��;���+U�S�s,�M��lؠ3�Z���s{�����R�r���ԑ)�� �j�2>����'sa�K<-z����9Fo�4��c�<�g���k��s�T��U�&�1��x�x�H[�)2A�b���
���!*���8u�+��x���Y��o�t/2�\!�_�V�X:���֣:.�����Y��ew����&�z�ws\8AK o'�<����&�����I�)2_٫+�����z��KЌ�F�T���z��[U�f(����w\>���":�B�
���'��s�T�yBn�'�z96�E�)�p�aq=,W�u~KS�2���V�D%{{Όfoqٌ&�(�=�%�Č�tg�� �������C���|-�/���BgNV�xخv<nm��)�%����뫳�k߼�����õ(��g��qH�+K
�s��w��.�{����^���4RP�lH���y����L\��N�7�h���Ȉ<�j�Æ�vXY���U��ss�Z���$�eѧ�dl@�*|��,h�H:��ܻ !��V�%gH�|�e�1���U=/�ޅ(�r�{�[w	ۈ�vI}-�^�k5{6�oa�Q܀���Ɲ�U7DH]�~5��'�B���܃����8R6�BgD&��x �)��=-f���Dg��N�\��	F'
�c��B 6� �Q^�,�W�g����c�1۷��qZ> ���W?�,|����(��Ԙ�U��z
�n{E#�wQ)F�/B2���؄��3-Z�?"T��^r���~bC	a�Y'�}�&w���gH�!�@�/�`���/�c�T�����P���wi�z�m"4�`�6X��㖀�0?ֳ '�u���N�!OI�o�ش��&�
a���ıe�'J�w	���đ�#����½����-��g���aЈ����q���[��^����?)�D�K����o�q �õ�`C9��`�A�>§T?�����l�A�TY�ڼ��D��.P��<3hvZT�\�;�[C��{��
���)�pB�o��A��7��o���~$G�@J��dE����z��5����a��̕���ԚP6>U�+�j�h���$���i�_��E.������g-ğ�"N������<���8O�6Q��`��k&�j�Vq0 ��:uf:5��^�m
��K�#�u�b�>��P/��+� C>��sn4���5ܨ�L����e�[�İ�p����Ĵ6�' ���/��{�A�->`9 �=�ۜ�w5�Se6�!ȫ{ ��H��w���R�=�%�\S\!!|Y{_��ġ�M%d&*��V��|�7>w������;x1[���v����nG�3�w7��
�j������kUr+�r33~��I���72R7q-��g=�#�'6��1��Z����s��in  ��s�s�z��W�@1Cf����DFW�?J���Y&����F�T����톙?��֥ۑ#Wi˕MZ����������<P>������sͰ[���GN����\X),.�?y�~]�:��L���n:+�-mLyԶoyyu�k�L��LJ��Zg򶵬��g"/D��3���*[�;[��K�g =��?=��ȸA�X'���N��}�d�� ���$��Jb٩�|~�L�i�¦v!��lw���׼}��-([�/:s;�\�@�}����_+�3��/ղ��Y�X���{}��s�x�D]{z�[�i"z�^xU�8�_�� �>?���F����XEPO4�&��i8D�s=9K>��阂��M#2��B��A�9��f�z������1f묡�ǿ��ތI׌PvZǥ���\X������ؽ��5���5�Дy�9���/J�5]�N���A�3�x�(.��G��"�ݔ�C������|�2Aqr���fK�����H��^�O#����m�E?��W����e�KK	���̗��8�J�Z��v���S��cP$��O���|Y�a���z̺�pu��3|Sei����]�̧-6��x�dcF�o!sqlY!���DE�	�Z�]"��	����qJ�����\g��ha$`�]�|c��qOXYh�H�ɒ[-���րf��Nw��n��p��Y��w~��͝ ����N/��_ P����"�]��������[��Q�zQW�ky�׀�[�F��u�
we�i�i���+k�ҳ��V���֔�2[�$۶�:�{]�k�.ƻ�5I�W���E�2y��t��l)ߙ��.A���^���kC��Z�m�6D$`�w��e�v�A���#7ɾ���<5 <�m�Q1]ei����5�IA4d�.���L�������m������P��a}Jd�V6e~s��yYn¦w���U�O��U5/�>Z��v ^��c��)�I��H$�P�,K�"+�~ִ�'���)Y���羋��k�o��~6�$l���
{v�����	�0���"�ճdBN�iĀi���)�G��̮iCCx:�ay�|š$����r�<\5�=k��*�
�	�Y^�BQM��Z��Ƕ2����jh-�<�f���qi�^��6��1�t��+�Ql{������L�W�8ta����ʼOm3]�:����,���Vz���Y\�Nݡ���T[ԇU�+J���6��u���;��(y)���H�ч�J�6m���B�g�9%B��g�"Oe�G[�,�ګ��	=v�������q<Q"���j8 �)�ޡ��=-��۰M����q+S�4���lV^jh3jX��T@�z(�9�,��r����q����_��-�
A��:�I��J����>��cz4�#5[L�z\�)��fYy ���.q�:	l�	���=��������L�5^����(h%7S��s������X��W�!�#�h���ݜ�� [��3���?6J��=�s
�Ko�$�-%�����﯏0�[��gy��'���i4�y�+���n&[`�A�-�=�����"��2�!�&�w�0dr�/��(��HS��H8?�c���P����b"�� �o[DU �q3#���w�|�X�^�u�k����w�M �X��R=D��Eϱ�ћ��n5�����w:
ߵ�-�)WW�_1�E���U��(JG�Z��v��X#�Y�%�^V�ș�ִ�eO��}�c���W�tam�������p���0��{���_Bzp\�o���Q ���ϐ���\7�@������\t��@����l������P�-A��VS���������Vy�
e_p�ߣm�
e���íiV��9Xlitu�4[�&Ҹ�2HvNd��XPYoM�OLL�e�#�Ȓ�'(�����y������E�";+�+�W�`��)A������N��1,�41>2*6W���N��q/voN�	��N���uzI^at��E$J���{��'b��^4�`O5��X��x��zPH!/�u�j����'��8n�ʍ�W^Է����ѱ"��q}�qXm"�Y����}X-��ݿ<FDYp��WI���cQ�X����������Q>"��J.�7]�C��:�+8I��<��% B2XL��KM�F�k�6��%����N�d{��yz�X��<V���\Lf���֩+wʫ)5��6k� ����%.���9��v�:T]B�7W[N��Cn��5)��U~�
�ڢ�IN�ļ����ew��_��k�Q��)��%��HÂHm���n�
Tc9 ��*�J�Z.��L�g<���Sa����Wv*!'g�Y��^�[�w�g,͠2-7��E��1��6�/Qqp8��y(�F�������^��,���A�#|_�թ!��.���<��$`C��=����3��S&��5��R!��=q�o�,�0�Ov�wRq9})�������㗔�&��Ӈܵ�^�|'��ŷk �_�K���|J�oO/���.wk;�Վ�|��i�@�%j���ߵQa}�L�!��Mת��>�2�f8�1�Q�Rh�%��@ꡤ�����.O�>�:��}]�4�d�#�� �$����[�L��a_��R�sӰ�xYlຍ���)��J=�s#
�b�H�n#r��5��y-���������v��p��WkG�����
B=��?���(^V5��Qo�s�G{�kh\.��� Ƚ���D��˪n�j�;'��+�y�T����o��e���+pja�����q�:�{ш��]>�#��vT]��\nx���֑PWu�)���*��hb���R"��Rʴ'b�)��1C3V@Ũ�&Wѭ��e3Wo����5�w���j��L@�Ή5��/��xV�(U���擎�)~��U��n��7c���t��=B�Ư9�~m��� Ќ۬`�ڝ�n鉢-3ɌG�w�s|�_�?S���SK����A+E0�b�'L�'{<�N��ΚL��iµ��%p�?�
:qĪ�FsV?Wʵ�P�A�(�"�� Џ�S��9��u��
�;���~}��Z�*���d�`�)NN��p�J������v1�e��t@�N_��M���*u�P�h� VaĈvAⳔ&UQ�=s���A���P˻�F�&�H�
�����W���N�����Oђ#{����us��:�,;Q�*m�6�$��2E ��Kf�E���}<nl$��{�}��NR��8'U�n�ԡ��wSX�>��Ъ���oG�63�?w} �b���CB�`��E��}�wM����B8gbX�L�	d��^.O3�&)��@��O��#��c��BΤ�Nh�,�,��Z�))Q���BM�'o�D��R
�3V�t�^���A��A򖻇�k����τ.�v�q.d�g��יL�����D[��/{��w[�&ڸ�˧���s�fr���{�����t継�}�زhR�˗�,�XR#L����� x	�9�$�MW�E	^p�<����s�ye�d*�ٳ���h
�4�zMWy�|�T�����q%vɷ���S�Un�o����6��v��]�@�i��a�ܶP�\��j@�ƴ��@��uP�m��l�?`ݣ:��lk�8�vH4���.�(u\/��Uk�^.rY�1o+������& }���&�p�a�"���3�bY鰮���:���W�Nx#��(ʁhv4��g��N�&*'Z`�^��o���	'+W��Y´h+�v��|�<I��NtǠ�=�B
4�G�A�n/?}�~a�ᤴ�bPa�B��*6�Q^���n}R�⿿��w (y=c�+��[��ay(�>)����R��v��d%99:�$~�����A�?���O�Y���؃����A�6�4�+I�zǢ�x�O@�s����\�N�r�)��i/Ό�Ts2e��V٣|[�c5m.��c��-�X��BM�iF=��ú���q�<Wwi�B� D�%8֖�;�\3إ=P�;�A����Iz��ndlq����2u�2&"f"�����M2n��y6�Ĺ_(�Ls���
�񣝣q�<r��ܖV`���!���G��ov�brh��ԈО;�>7}Nj���0d X���&"*ܣ(O���I��ߢ~
{_�ѓ(�I*5�d���I�c:2c�_�o@F�iO^�*�y��?�����]�N�ڃ�׺dn�Y�
�X��{ɰJ������{f�W��ge�z0P<� �[���RQU !'��L��UX�@d��Q�ѣ�R���y��jk+wV��t0�-i�0	>z7�9.�S�#}�N���j_ �kq�C�l���z��U�$�YQ���Z�f����m��	�)���%2����u٠�漃�\�FY7�P*[�Խ���Y����#I�� �q��KmN��0E�)���L�LQ�k#}�$��N� �'��_WT�Cz'����!�k?������y���� ��r��v��Vj�N�
�wF���t��N�7حO�k��,i���&��b��Ǩ��qG���5h~�o��G����'Z�'�ӓ����#���c����=�Y�Z#>'w!`��f�3�v7Ì&e�f���1��Kt>\�Ǭ&����'���-��5m�£�hQ�2qb���'6����]�q`_'"�"�<6F��kgF��ٟ���C{�[�T�Uj�^���|`�E�
�#ES��J���⾁i?�]�J#w@B����'ʾ�V"����X$�}��(\+�d�SI�3	���(��ȱv�h��y� 'a���g�n�{���+e�'������If�O(
P��c慡z�u���>�����Q�n���I3s�|'�e�k�����e���u�8���g�+h���+N�!�X@݌�?�sS��|Eq��/�^s�<�c���G'�Si�)��b5����ן��症s�q�Y�"��$֖�̉�y乍����?��_)6<�b���4�3v���b�2w���e��P�tvx��_ Sr�p�e�
���6������}R��ɲ���1�Nۛp}�tI]�4�ew�2�4�5�V_��?�r�&���Œ�s�S%_�NE�k�+f�7��<^�l���u<@*�}�K(�C��u�
�iz�?~ �O/�S�w�K�����P����Dx!9��g�J*g?�M��`��+R��x(a�^��C��sv�(o���~ܨC���2ᷔ�TM:��j`tᱲf�� }��M���&j,�/>�RJ�mS_�{�;��.�]���&v�>���ut'���
�q�+����v>���i�7!���g�9rK��#�q�ܚ�{����-|z�~��?��<���1�Z¨ 9wO�p
�礍0�y|��V���#-_��4s�t���H�MQJ��ܜ�'B�zX����-~.� �8��M�r�@��>�߱�tT��YQź85y��5�^�M�ą;�9Yl�'���Y���������XH��0 �vp�A�g*Z�K�k>�f��T4�l���v�yq��(;�pYXȉ�� T,.�������0\\C}g5�՗0^�1��ȣ�/fc�n�q_��f��R�T̖�1y��8�wM	�8�8mt�8{�,�D�v�1N�-���[A�8���d��D�ܕ�M�t��F@�~�[cZ��0�)$����xK~9�B���s��#+�`�njr�=�A����Io��
˴yE���ka��7M?�&�]�`�W��"ǭ��N�:�pQP�]64 �D �i���wv0b��iglU^oY��Q;��8M<�>V�5O�U�&���wt�P�5B7*-Ջ
�7v$����(à�K����8n/�rcq�]��}1z�W�<g���5$��D�d�#��-A�QCc4Ix��Y�v?������d��_dw�V8���ҏ�S�.�d;��1JW�m���O��Qޥ���K��0�sѷ^����@��Q��и�3�ǳ�S<(HBG��p)P���!�$�#�A`qݞ���*��I�d"��8a"������[�C���P�"0xk���'8e0]z<��v�a��d!��J�I��>���XY�v���o��X��ڣ�����5&R��4y��Q`�[��&߂�)*�Ro3�����WM�6�W����cJ ;a	!=���Eڱ�6�S8sIFߠd���z��}؎��L�Ny����b7���k^ם螚����e�LA�Iغ�5R�@�O  ��� � �h��%�)�N3z�a�c`�m%�\���YF��2�ӟ��Ξ5���ò6�Iڒɕz؉*�cAu�؜��E���y��Q��f�+��� �Ʉ9�J�PUuZ��{h�š"�
yM؊�g�<xHe�#@S�V'�-� ؍Ň�@ʹ��p�Vb���!0]�KzX�ē��@0�Z�4�6N�Rl����ʻ�B���o���xd� �v@̸�:�PHb,��^h�9O�`1-�����N�dv��=��V&úKzu��!�d��ߺ-��IN�5�I:#�L��q�}ly�gc�+Y"�����D�z��7��Y�B��j�`i�����{p'x�@�M�n�7#�,�\���G<-TC�\cZ�ނŌӛLd���}C�Ju������c9Bjf8��c���7Õ�z�.�
3#���ǓlE&zwۑ�:���� �l���WK�w3�x�]N���.`.����IzS���y�|�x_�h���7z�6��3kw�=R4��5����]I7]���:���l����k?3hE�&6�Z�+ϼ�;�\*����ϼi�FV��p�����Y�ʍ�^�+��Vߪ���Y����P��3��]Xw_a��h`�|������k:ڒ�Ҕ�0�j9�~����9;��Ӎ�PGt�E}Cn"������6�� ��h�dwmF�/��$�y}Tom.�槂��ߔM⯰�� z��H���oE33��G�UN���i?�s����.�jd���a�u�~O��~���z����X�N�Bs�ҞR`oY������5���>�TD��
0�XV��J��L>���6�8e]�B59��  Iw�"�iN��mNX�óȉ�j�t�\ �%�)�Pb<�Ȃ�L����	 ¬F�[9�(����Q�K�%cb�������9����@Yƽ��c$ޚgJ�R��������~O�M���؛�qC��Q�B\Ѯ�lt��W�x\{[��^��M�0CS�^`�hnGf��8�-��_�V�����=����|Xv�o���hy�m^$�1YE ��y��>��fy�r���e����~�%]d�
Z�l��v%��s�k4b�0G�&H
�������E��_-�l�Sd�
��UV��3F�S^U-B�^�oѴ��u���y��3���Ǣ1�(Զ��r,��8�0Sj��_mm�p	���j֓}`=���B&�`(a������qoO�_�:�WY��f1���qb��~��Smp-��r_S���B�5�9;:~
�����T��eQ��_ZB��:?:l������XH=鷳��-l� +���!�Y�W#��B;Zt���i`·f	��+e�N�B�s-����By���f�VI���J}]��M�*^X�ٔ���z���6ϫC%b�����}����wEb����;I��Sz�e��L�!"'~1���6�v�W���]�Y�uȷOCƪN)����I+�,�Y$�R��;gv�Ȧ��Ue�a]�f	�_mJAG�N�X��<�C&�T�����-,�zX�Fe}}[��9���� =Y0+5�%%�q2	�1�_�x����=�<��#*i�)�DTmg�-�e3��r������U�C{��^�ڴ4��ө4Ä�l�D4`ea���@8��*p�)�v
�3�Ρfu8�=6�p}8$&9B�S\"�v�FSޛ/��+PJ���*��\L��EK �sdB��}�lf���Pp2�����SՇ^:0p^�"��ib�^�'A "]Z����M�����Ү��(SV�W:�ѹe��n6��ǁo�c� ��y��x��-8DG���b�\;_�r��ޭ40��^�;�(����n{��:���`�A�I��(h����	,�#�O�_6LH8� V��`Z��Uk��{����r��br�ּ�%�G�~6�������i�B��m5?�I�-���q����B\�N��6y?Lo*���,�劐�^�׵e˭*x�}5]
�����ж���Sj�b�#�����mE��v��4%��opS��s�8�p1nkutA�*qi��2n&�9: eƝTr8��w����2�lÉ��Rl�����$�PЖĻȳv9�{b����g���_����Z��8�q�+�FH⹥���=*��ļc�.�0��)���x_ /�X_ԧ� ��0�'&�*���U;�}C��(�F�ÚJ�}/BtN�dC���~�����ʹ׆fH!
�hr��hW-�ń�<�(�5>׃́�G��A����P)�M�a��DS�]>D#A�Eΰ������o�7{̀�h�f�$�����"��OB��	�Ӽ�ټ9����`���#F������C6bn\�ߩ��U8�IL+��,w`s���*��p� ����*�ͥGOt�E��Ѹ��A�ifC��a{�o��;onCV������`t��0?ЙB���](j5Ǚl��ͱ���Z�
�C���O��Acx��K[e�e[\������Ux�/��]\���LyQd����lΫ#��EFk�f�ҁ�ۤ��2:S�$u'��T�t��ҩ���|t�a5^�E�/�8�-Vl�Q���h>�w+��RΟ�,�T嚡
�g����(��z�!Kd}���7mJ�9��n�~�5�o�MK^ �%�}S��bM,�~ŌU����/�&`Q}��^[�k��O���!w( x���X1nT&�Q�����a���_^
����s�<���e�hS�<���X���\ދju�����#�ڬ�Ľ'8���w�����J��֘%G6=�ܹ5�2�h��Z۸e�+�HWJG3�r����Y�Ss�����^�������z��f;�}|���Y��w��έS��Xu�B�4���1OjKq���C^f�q����y�����l$̤�!8[r�K��PU���O����V���~��3}�V������p#k|nB�[	�^���"{®���m��4߉�fv/Y�^����]5�1홃jI!�����b��Kv
�+�ؤ��Ïr#���z��˪;G�M9@��S2��ݘ;����i�0�݌OK�&��mq[�R$�^i�� �m��m�g�}�N����ٵ8�$x�b%-͓�w���Hb�O�ez��!�4L t�,	�}޳�*�ş\���u�R�`W��3-��L��b	!n��H�8'��n��S	R��C}��`M2k�[�_���z� ��u���餢�h�5����tA��qu�x��*ҟ�:���yt��A�A���͈�8ζlHM�cVh�?��%�L��@�xЕ����ĬK�w/ݜ�H�������L���
HR!�����ayM#���}�x��{�r�S=�&4n�̠�V��B��p��Q��������#ھ��²� {�@�/6�o�X1������9�J,dh�{�WMѽ�99w�ޢ�ƒk�'ߦ�9wն���e���y�׽F&ao��ăE̢LM�xV�"dW�J����V���K�Χ�^j|Yw���Awu�譓x"<ǻr������]�iԐg5��6-Z7�b�|8ﯰ�N��T�^}�b�E��%߰���*�}�뙬�PW_Pg�wftp e�"�TC$��k��O��pݘ��Y�����h�9*� d%�q��}w<�k\�t�wF]��)p�����փL�}]i����S��)�/�� [<�E`���7�a`i�u��ǂ8�ܶf+��rr�u�ˠ־�� �ɼ	}j���\F��^w`軫���m�")S��9����!f������=�WgP+;�`�!> ����ɳ����K�����K�� K>��a��ɜ�R������eu!L
�H�i��m�#[�i)omy����梀e�)dGM�wQLzC�9)���^&���O��H�2���]d���+6'(>��
���ReA�oO����ZK
w&���7�<�x���(� ͉������O����:���^s(�>�y�A�m�r��@��t�wW�7�Z� �Pm��u�Aď��J�{��n����/���o�!�_Pg���8�osƯ+d�5n_<�����d�h��
RTX�rK�|�[n�����~��'��M��o4]n�e� �#���;SxkĆ��>�̈˯[�B�SL��K�.�_X�Ȍ!i�w4��_��8Cs���c����n��A�	҅�do
A��ܜ�Jp<��;�pd8��i|��a�����W�j���\�0}��0�;*
]w�"�1Zx����+K87wÀ��``�$�6�?$؀���%��d�=��@%J��E�y�f���8��Gm��W�;{\ZEE&���`�5�����Hq-�M�[�{��慄�	0�pC�&��Wh���%���('���.+�?
�?g���M���R���e)��;���e��툺�!Z�7�
;1��k�C:!A1^C������٠Ti����:UY#�>S)����]��uU-j
ݠ�kV��$�.������C�W怟>�z�	���<�Ef��$�Ⳟ��#�>���a���\�cp�u�х��T��%�z sE�&@��4�/¼�r�y�m\*�yu@��~�l�qe���=%���9�6 �y0��8��������Y(���asD.��/a�9�ݏ�Ѿ�z�'����uHa��Z�j��'J���>�Ng�R��	V�t����%���%�#��j�B���[��k���墋d��jdb���=���W�њ����?��ϊ���g����PU����D�T��lN"j����E$I������S�l2�Hzi�/7�Ju����cϟ��S����1A���O�U���f r$���J��{����%U���07�m�C<|/c]�U�ܡO�f�s~-�	u�a.}5E)UWj�´}-;��-`)�ȘEh4k�u�r��?�'��'����?�F�pt![H3y�H�Y�-�X��{Q�n�*Ut���ဒ��
^&i�y�V�?T��P�[�S�W���,U"OĎ����ߞւ<
� .�&t�ɲ7fx�Qa�0��f�;��62����׭_��̛BQ�~�W���4��6�Ti0�^Y��.p=f��������LdD�7�w7L��t6��l��>��=������1�\�
��a�w��~3h����	�4v�G��N;�B��G�[Y67%�s�����aH���)���@His�*���&(����+�~����?%pGri��D:B�����]�O)ˬ�r���ѱv��)�i���8ECciC�CQ#�ow�73Sa�. }7z�9���)�HiA�}֠ �ˇ�^�+4y�q��ѩn��5�����wE��l������a/<sW�[���������t�w�1�(��'�a���+h�.NU�m�e'X��rL��?��t0?j���+;Y`��	v��HM@�p�5HZ��G�Y���i7�c�H�lY������i�+���� �� +^��p�״�Y�<{u1��ߑj�Zl����q'T���Y	E�����-����uS^�W���w:���1S�	�L��v7J@i�7��W+�D��kBRѶ�yh>q#汁a�v5��u�P�|�ʜ`͜��s�x�.���������<,�Y���&��3������	�x]�?~���<�� ��i�W��u��;�V�M��M�5C�[��D�x��i�*�Ӭ���k�8*��nO�>?�|����FRr�}�ʘ���϶�7g����S�^�F���4�{��߀��()�]��Lg��ęLk@��X,�.ٵ�ۙ�-I����=��h�����{��l@{ͩrʮR񢑮�d7˵�O!P񢀟�8ڴ��F��M\�[�H������Cز�eL�����ޚ0Qw��>�T��O3;��=�о^G�a��oҋQQ�2%�#*��eK��|x��:SBh�2w���A��^Q�BJC�a�me�}DrV�uS�M��F�M]��v�P(�>�b疿&��U˸�������ᔰLӔ��� _��{��R�:X�o���D��iP���E�,7b���Wu�TLZ�'�e�������[3 ?���6�md���H<�j͙`�B�԰'�z8��ʸ|@TT��Fg�.�����;Y2!ī�-gH	hs��V��tˇ$ԇ�!D��}��ɟ VETT'�ԟ9ʑ�4���|tD䜾)���rEGi�6(f�L^	�V�����PY;��
4�iV�����[�Q�o��,,�.ܫ�l�<9ct򭟎2�0����afG��DЄ�&I��=�XxtlAZ�T�����!�+�6�P�5�D�٥�;�y���(��{}�ѭ����9.Y���}��Eʼ1�J�vfЈ�|<Z���cY�Q۳�«x�<O�%�s��+a7�[���I��������G:Z�v��1,��ԫ���PU��c�o�3�w]V�qC�i&�[KH���Wx�������.k;^�hd%P�~V��8|�@�2���֋��J�����'�|��������-���-P�'��|a����x#��Y�ƅ$�,�B-\����j�ET!mx�8>��[j�mVʎ_��2B�ξ�Z[T�����h��#�_��*�u�ԏy_����9�>��e=�꫻������U��>�N0u��A�J~���������$�7cZ܌gG%��_�9��z}���p�^ݟiW@����k��ܷ>
��#qF�K(��_�-Q^���֘蝌�[�����e���n7睊���� ����C���Ǣ����	����D��	�6���c�u�㳧���{�/���4<Ҝ��f���@Gv�<�)׽G�lX�J�m�Ǯ���;�T2�;8�aJ�3��،��e�rz;m�O4��;��\���(U �=�-}P�$ƵY��g��Iu��h�`�4������V/���dd)/Yˮ�^��fG)�
*��4X�Xs�ۻL�;[�0q&���n1��iX�i����y?VJ6��$e�o��oH�l����L�=����|�x���.+]_�M�?2�'�d��y���h��| ����c��87���k����mVؘ�S�>�І�n���V������qAnP\��ܹ	�sy�0�τg�'���v����wu�3O��_p)��TZ�qܝ�KXR��l���݉eyV�_X�
[��R���ަ�GNh�{��I�	�|aD7�c �n#��r��? �Rʆ�Y��
"��O�6!�*x'���^�6G�W�6&3/f8�el���nv��Qk�Gk�"��Ǳ�c�F����7.�_���]�����ɾKU�n5�H�%�-�fw��J{!�(��
 "$�~ؠm[��ۿW���
#	K/�{��KF�n��%].��zF��`k���\Z�P������tA1X�-6����}8(.�$�_kw�����S��XW�����C-%��t�V,�g`?���3�ls�*O�&�V��k�qT1OSX����D#��d�x;�2���/����ZZ$mi����"��6|F �ı��0e	f�@�X:�Ż�5��cp3�\��&�N�w}��*?8�)`ܸ{���)����&W�)R���7னH����ޒcA��Iu)u9a�۾��o�F��{B�
�ϗ�+�#2�`~ײ�~��6^��!�>Om`9t�MI�,9�JKy��텚^��g��11@?`@C���u��A��h�r!�x��{������(4A��o���Jp���Qou"��ag7 �v��,xG'��=g��1�O$91�6��71��}��s�ԛ�A5>N�O2H�
)Q�qtQD�x�fX�:����s��$K��ܫ*�y \��(t����M���Ē������y�q�E�W�.�=(*B��2��2��]�t9��_4���oǍ(��Z����N�� l�O�c	b�I2�Gl@oG|���K��<4{�t�f�wdBI�y��l�?j� �'G�R��{�p0�s�Xh�ugm�O7�Up����Y �˦�pNU�$c��RN��^����
�zF��uD��Za�<��d?���i�鱳��r��2r� �wO"(��f�p]t�%���l��}�B��{����+wFf2����o�ocu�lA�Cz�W"����j%���U^��������lEV��<h�ćz�S�h Ɠ�X���T���n
,��Y���As�o��#�h(N�˒]�
�8�OJ��؋�Cz�!m#Լ��O�/��\s��Q4��M�(�?��V:֮l�qU�j��W���Y}��wY�3���T���[c������'h�a�������]"$I��P%t�"?��G��r8���/�G�B=;��\n�;PϐeI�Y���W�Ud����C&�CZ�´�
�_Wf��un��� ���z+�B�Jr__���G�J&M��i�' ��%L�P�%f?(��] 9�Z�<�ش��D��ϼ������K�3���nN���p�D}JNzcr��(��y��Y�%���;���ݱu��ح+A(U�����4������\�Q�v�^��f��ހ~d�q]0l ]��C�n��1:��2��I3_�Tx#P��jflA�Ů��u`9�؀����г�*VN�\J-�����G]��A>E���K�5)þ�H	; /�'`2�����ML�,��9��W�J7'm���K�D��eV�� ,y���l��&�
�bg��2{�����vd��Q��c�=��"����g�~��9��鋾��WA_Q�e)Ѯ�{mD���Y�/mznhk�{[Bo�?�}xl����F}�/�["���)�!�d�C94R��f�G5�*��jXn3)��M�d�2��I^H\�6y����eq
����� ���x��=��fu��D{O���P��a��E�ǳ ���B��'���H�c��lt?n*|j�I�p�2I]&�@B����8��x�QU`��J��ӵ�P߶|/h$w�5����9�Z9L�P���k��<�O�AC��B��h�-<��-�%r����F���� �#[�j��a�*O#?^?���[�;ac�P�t�,�V`��=���w/<oԗj^�k-Ou��r��T�Xٵ�cH���/�}cþ�`4���C�-�@�^_R0�.e���wSs���e�Ru�,��1�nnc�{oGq������h������h��8~�K�`|�m�ǟ��4�$�3q�#91�M�]%n� K$���-x��w��=�5ZS��h8��O�ٗ��Y�6'�vʱD�bz#�KU��}\H�*R�;�6]���^���Q'+ЭXF��l���Wδ�i"�I�5u��à`3�P��1�t"z'�)���y���2�rѫ�A�(vJ���;���o�"MZ�]�o,g����VkT�瓄~=�9u,���ձ����s�Ɲj�K��e��)�)Og�W�_�wË(Q�0������T�*E4��U���ɏ�6�wIU���~(['�j,jl�nB�B̂�/�o��vp��>)}�D{ZI�ƌ��M?�;�u��쏗!<�\���u�M����$ ���q��