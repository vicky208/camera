��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V�h?�xrMIp*/�p�x�'�e^~��?u�ik(���4p�Pݐ��o��d�m,������i��p��1���M�f_���cK/�Ʉ���;fGz�2�ԩCA�4�ŵ2�{س�
"y������U��<ÍJIA��v%�����d�9p��'1N����\�����t����eAI����U�\" ��`�@kD��<���}�9�2�pyK�뫐�N�yE]� ����K4��M��V-?)5<	�I�Q��xuq2�9�Yj�g��Ӹ?+�Uvt��?�Ul	�s�r�e�`��E�)n�=����]���".TM1i�軩?J�[����؏�yI� Mn%-�� <v�t��]%2��D=뺩��̦�#� p����)��\���BK���Z�bZe?q��&�LOlcm�\%��/k��+����Pb��D��f��b����_h�LG�/0��ٌ��9^*gj�X�d�;F;HJ�Y1�S��ՒȢ�w���p�.����EY�J�����J4�7aG�j��l�Fv���'�;^9�1��]�I��1��K}Y��)���3�K��}$��]��Q�4
R��*�Ձ��ё���k��,Q3G�{kQ��g"��9=� �=���CoBwt�3E��z̑����Ğ̟=ӯ!��|�J�'C���(���~uA��Uv���ю�P��졬I�&�`�u�,�-��K�u��y�
�k>T�Y��s��h|F%4O��t#ڋ�؉��#����-�CG�<��|���M�S8�:Z��L:S������ ˮ�+�r��$7�W��ߎ�'~@̼���|���S_p�N �)aje0gޯ�_�4�P�!Y�'{_g��=X?�߸�n㨎�_���A]օ�����|G�슠�����)��S3�>��_ny�u�#Ͽ۔�(ɼ�2S)<��60�A�
�E��J�W�@tF���ځ Z¢��J6�	Ȥ�3������I�%(qZ0SB�1旃8u�C�A�葧�1�;�t��3�J�y�k^�.�G�>!q~���c~G>:�A��@�LT�X�r�2��ׯj킋�R�E� JP�����V	�aK<�ֵ9���⭨6�*v�hzT�%�R��s
�Zb�s��JdT#�ZmۅU�a�v�v�[.�����'Hd��H�*Vĩ�Ef�ù����E�Z58��U���; ��L���O�r`/�1���m�Ψ�ż���}˘�������U�F�����O��8>Z�7(�̂r�g��v��p��WUY�󞪈�9ץ�b�始�AZϵ��<�\E�!s���.	�цm��k�N״��!�)D���!<�y�>�ؤ!+�Y�&��j����Yy!�)���Iӊ6��܍�͐A<`�/E�c�^ޜҟ��q�AǤ�8���j٥U*��㰴eOF/^�o�n(I�$���֐���3w�]-�H-���Y�+R��TJ�I/��{]��Zv,�W�97e��$����=o}�Js�p-�	+z�!��9㬻_�[�\2�x�cF��0�ur��������^�\ƇHj1[g�C��`�#'5!^���(I85*�_�u���K{�(�o�q=��`<Y� ,2�徚{S�Xԙ��L�㡇s<�N3X��+r�[�L�����
����ӍZJ���|��������^yCNԖ��KP��xq���4B{D�=iGX5�Z�)�:�X+�S<��x�UdC���L�TeV�8������KP�ls�����䮖Da��4
�N�nˢ��z�C)��'�?fA9��I�0��1��8~����j2˚�ҰA/ߣr���^b��Qt��R����,weq�š R�#�`Y�U@�LT=�ִ�L��圿��iM�X����ys�qk	�c��&!�o@����������!��!�Rl����׀�:�&���MJ�<�3�^�]P��"����_��-O����T�x���K���poR���<�f3�U�Ond�?l�2���b��Z\5C���+�u�TÊDC#4D�;���W��9�{�p���{o�
�M��Z���GK��Pt���uHR��9 �C�N�S��?>yZ
K�az��U�bb� �;4�=$, �Y��Wa�a*.S�9��׋�$�Lx	UT���e���\���|���YB�t��c�Gi�3��0q),���� �&�hD� �eۺ��?��T�!W��-��0��
B&�k̻�"K�G��G��$ؖiaM89R��c��g^uo���s�~�/u��9z�Q� ������U�f������-�v��ι���ؖ�x�]6��S]>�֯�
���w4,�����&Y�t�`�?�v*���h2m����é(/�h���M�7im��9�f^��xv<i�Iݡ���G¸���ġ�jh�����R�R���>���z�QYN:���U�1�/X�H�������R�|�����H�he!78`-):J�H������<i��Q�꧐��ꡋ[q+��g�R��v0�/˺�潼�9A�Bo��<�Ѿ(��k���6~{�ف���:�4D��[���e�ʡ�Me�*ꈲ�@P�m~���U��w�6j��
��0T�k�Dh�����f>�6M�\Y�i쬢٣UV}��Vm�c�3�hvK$X5P/RE9g)��
��	:��S�1�d��1o�����8�ͦ�+I a���z��N�5t
�;�M7�>�v��Hvff�QަcyRI�Ӥ�!�Q�G����rnB%�ẚRA ��1�� �4���0��~�	��u9�{�pۍ���Ȍh�&ȳ�aA{��M5��]���]�{��������T���t�k�ߺ��+��I��Ǐ�5���l����הw�ǽ�L��]��T"�r03%z�KFNȐ����|-��v:��P�J�m�W�a�i�r"��� �L��<��7*k9��f�ڇ>��{�1���.�D��͈vi��xԉ�k��#s7 b��v�/�y����WntT��f����k��7Qi�͚��d��eL�[�58�>�8,�Ҩ�فO�F�t Z��L�hV��tJ6�|�<��t������ E����#;ߙ�������-v�(��k�FB�.Ot�TJ�@��(������IdD$X�w��wF�)ݜ��cl���y�����͓�q@y�7��J[�*�0[�O�J�S#���L;�)�R�����@`�
�l�h�0�b`� 41��>�A��_q~IR%��P�\�K�5 �P�ۃ�^��-q�
��_�uz����Q�ms�Ӌѣ��1�o�EG���G�k#��Z�� �@ ��k���H%�ے�%k�_��4&�<K|�q�D�\�4H>��>�n���.�y��}�Ȏ���� �2	�ל�z3�O�>_�|���g��E���2ug���>�y��c��3��I�:�l;p� "� �-�X�ǃ����=Y���/�ji6?KM6��ɗE^a�4��d����f�?�Ѻ��W�!^�Ly`�pK<�d��~�kN����c*������R��u���(���FZx;���ᙬT��q����8���S�v�n�Ni��:Uxp#�7˼���%_���>���6\�VU\�7c�d�(�4� I*vj`U�G= e �����zf-9�\@^���x��*C����p�΋֗��ڡ>��ӻ���޹� g��)�c�{?�����N��IɉCL��K�8�}֊�����F� gx����A��T�������<렴?lXv*�?�(LA�����9�J^~�y4�VN��sR;����A�'��*��e'x�'%g��vA�*���8�w�%� �;9_�B�T�\�� �ߐ���Nъ�����*��Պ�cJ^x����K����yzL���6�P��L3�g,hJ�� 
$��]�	�I��cb������_Q�g�I4�-M���دW]y�ڂK��*�]yB�eO�`b��}�eW���W�ӈR�����=��d��S���|7*\	j�!����Mh.�x4qk-��th��7X�s`��XH]*��n�d���}��C�s��Ǽ_�a�R$5=S��/�=K[op`��5d�6���ӈ>Ց��'�'�0'�?+�bK�׺�0��H���SNl:� ��57�����
�m�+[�KȰ�a��뭫�c�f���1���sY��A��H��)^��)&N��9h9aCU��+�$Ma����o��)���k�U�v��82�s8ҤɌ���[O!�j�H����hȑ��[�ۮ-(� ���Wb+c��U�e�Ay���G�m��֑.(}�����F~ȜN��B�^������)����h���|����Ik3���n	QZ*W'˪�6G��9{��t��!bf��z�Œ�:�;⊘�	kṐ^݈�C��KTv�`�1��&�������Ş8�*�̖Gv��dM�p,cȝ�
;ӁGe抩��Q��B��/�x�0��ڇ`~*'s�D1k7ȭð��y�9��/S��˨Hb$�ĭ<jg��������'
�Ϫ�7$����������_O�fM";뿊�F�z��Fl,]�4�y$�e�˴Us���	�A�+.jl8&�ݯ�cf��IȌ� *O�<%h?L�����~~c<��ݶQ��p�D�j����� ��f��k�Dp�h�t_3O5-)�Ҵ�t�gGZZ��fC�ʫ��C"���,*A�:1�1��X��,�#��Wk}P��8'T�n�<J�WR���c�^��[�ʪS�d���9meS�2 ����ҁ���"��kߖ�.m��I�r�zL
s`�ذ���yZ@I���H���5�a��B��G�_�Ћ�[�J��0��$���k�`l6Ò����OPf�b�O���6���g���,�o,����+`ԕb(Jh�@�Οc��vg��t�A����A)��ZT�&�����+>&)Z4�D���{ח�I��@�l<x=���W�݇y`�j�%�?ji�e���S���i�1ܺ%�>�&P�Buݹl�^Wβ\��)��X^dB�[u������Y�r�푣cN�5��������0���KU�f�m�T�7лZ�� I�K8�����x��s��لUҝe�4Ky��.lB�}6
�E?���a�ri��B8��gMmE,�����p�lP�3<�wnN�J.�%��zL��*����+�D�dA�+VA��e�pDOhE�l:�=�F��Q2qn+�%9=g	}>ӹ�8��QC:-
�-�w�b=R�8!�,Kƌ��uݲ0v�U
%4
����nOk�Zoli��[�ECԑN�ۧwz�
�1\dcM�%�^F�{=�C�6�7��O�ո2�:�͗A�JZ�Ц�0�ÁM�c��n�P��"[�%������ ���p��Ͽ�P�<\`�w౴�I��F��ҿ!��s743Wj�T~�ۅ��LGf�Z�Bq���,�<�Ԋ�m;V2<�Z?��F�k��������<@t�vA�|ZD��3嶫я#8�`��pWDM��w��482�q�:���7��=)�/���|nmt�oGI!�ɕNm������iP��x�ƍN���W:8��A(F�k[���d�%��"f���Q�9��A?d��<�M/5Ҽ�e��%���`���(���A7��W��4MK��ؕE2/#5�t�l�y{���u�"�Jcl�����>������e&�`)(l�r���A�َ3�,ܩA�6�2lp."�������&��%k6ܪ�-�
cX�?��x�Z����,�N�x�MQ�4���~�Pz���� od�ӝ���
Ow2���*$�Q����]^xv{�˭����D�td���t�(�m��rՂ�0�����·Rφ�N���T�[J�u�zG�������{)��o���܋��p������aj�@�N4���N�=ʕ�8�����#D���SI>����;Z�g�t]ii�#f�ǌ	�K��ds�I�������Yз��l��[�z�S�[t���������N_��<�p�~�'��������z�e �zXa�<~��7����q�l���^�:\��c�}p4l7<}���n�G�g�OX�O<z�{/���#��H1D��V�Y��ޙ���	�T�1�K��?�L#V�)!�e8�J���"�;{�/O�D�[g� q�p�����(�'�v���9a?^�ux(�kzS^�`�;�����lt��J�e��_��7���2�B�B��@s�/=�~�Y�����SJ0�aw�Z5��ֿ�]���b����$j��r
���{RP�6n@*������iT�&eP��̫����޹����!����ĞMMd4/����a�޴$(�%�@v�"\����+(\���=k[�b������ld=�����q�8�j4�o��$PO���}��颍���#2Fe`-�
�)�*�Q�L�3L���k�r�^��m�l�t�o����j@����L�Cs�.N����dnf�w�>T��t�6b���b���5��C��Y�e�T]
;��\�9�75��,���n�oD��SĢ�G���M1*�p�	����5�Ώo<A^�b�}�#J�WӤ��5�(\�.* ׀M3HP�B�+��'-B����(�97�W+�"�F^�?JC�4�P&X
*�53�QF�}"��E�mL��>��pZ��^�S��w�)���*�X/eD�g|$f�����I��;5�����md���z��a���d+R�me�o���0M�W��_�g����L����5�|%R�Z�6N���y����%0Bl�Yd�'��Ͻ��(=x�V��J�{*�Q̘E���~�7�KǑ	�\��fH:.a6YA!V�8�]�#�i<�k�hՂ���_�Fqw�O?�<�vfae!�;��&���:��ڹ� ;m7ЅіN;O��T�V� ~ ų(��\G���sH�Lҳ�b�[�R:�(�G��h�f9��̒0�f��Ǟ��[���\.<�G}~+Ѯ"�y?7����l��c/��ˀE��m�dr�V=�(�z�N	>rZ���d�=�_�=Lr�*��r\g�P��,g�$��̊P�0Oϼ����� r�h�!�s0Y�q�>�r-�m���K��F뀮��wf`���v��q)�Wf��*M$2!�
lr�72�{g<䔱���H�H�}���Ug7��\g�~���?�����V�1��th>E��:%P�i�R��Q=�]�`ӹ��y���(�;Z����/)z�fSήYK����a�nWC���d*����S�f�c,ȉ�B-�_��^Io�QHS�։ (��j7�mv�}L�_<�sM��"^[ D]��@6��V#�@�zt�D�A��d>)g����(3���i���qN�T��Xúp"a�ω�2]�a��R�6N��iN3݂l;���*��4��dS+6uv[�W�̉���%Kʱ/�ޜ�Q���b�:��M ��+/��&16%tA=1�~�(�� TٌbP�� �#�g�x�d ğ[���Y�(`��� Ta 7�Iq��Sg�.M�lcRa�,��zD��Ǻ~?�)^�d�o��[}��Wz��1X:�p��yu�@8�o ���f��T}�(��[�0�K��TLT��C9Ɣ�D�`�;a��Bll���+���6�Q�ǝL:�E)�0Y��������Y�#��l�zb+�+E ��mVIf� �Xr�&���ւ�OL-�!����A�x�Yk��҃S�;.�P�vݦ�GK��^�����Y������4e��(�@��q�"��j���*���%���A�z�08H
��ǅ��\�w�h���Ւ��

/,��I<A��)��ꙩ�F����DB�c��@��{��P���M�u��W �{#
百���5�n� �D�n��r���bT�,���/Aa���%��vR{0��sc�|�*7N���>��Œd�PfC�Qy�}:�������0T�B���W@ ���^i�VvD�<���QT5�
���'�h%-O3W~`���P����3�ӱms���k1��B'\��[�d�<�K#j�,�9�^,��R���"R���D�:=Q���b��apK��{U<�٫���i4[j$�A�$'`�"q�.͊�����R�R+_}��"e7@G)V\3�W�e���	��f5���@�����P�g������;�%�|9�8ˍ�,5Δס� ��苌/B����J��H��V8��x�,�nt a�����Xz�y��Km����79�0��?��DT
e�}��|�N�ܟ&u?�VrY��d�ɹFwN>���>����͐�5���R��1rF�#��ƾ�P@��	K��9�S�8)(Z�rB��o.>BVI�'K�N��t|�G�Vf��K�b^�JY��
�F\#�O&��B��.ę(�V\�g�dA�<O�nor�R��ޯ"��2��)������8�bV�jpx�L74�;�gx�t|D�i�k����X���(����E�Fr�\T������tRU���99a�{/�y�Izr�Lє5��2_����?��>��uL�����'��;W<�I��m���Tt��h�Pl�A"���H�n�pEQU��G ��w��O�� Jγh���B���� ``z��XA\��a�,���k�Tت�E�i#��P�y�gOª$��)6B+$-��� �Y�R:&�r�Zq|o���yumQm#��O�x�HF�k��d[R"�40dS-hD�p��}����:4k@#8Nb��J������O�̇�������,C�-ۈ�\Ӿ��KR/Q<�^�1�?{!�=U~q���~��Y3�$��=���	�B�r��rҺ铀�Ź~$J��q�a$�P|T����v���~�j}����
b�|Y�ӕ+�|ql���V�`��Њ�5Q��2�*���^�2��W�0�@�r���(���ֶI��Br]�$G��u)T�6x��.eY�xeu��e�YS9	*0�f�}��d�H�!E�Sf�.��;��XxF��B�<�hQ�u����4:e�5��-�RZp�����2mAz�7�F�m�I�M8���g�6�)f�X�ie��"����3@<���rLyR	XdAB�1��Z2��?�8��;�3Z�B�	.41\hC��$�r[�ѭ�͔�)�`�r�2�ȋYp�-�^�����$|�CN��e�u4�d��U�ǴV
���GP��n;�cg�Z�2L�6h�^Fh�)
��Br	6۪ү݆V��R�RǞ��ol���[�*W)/$Ys��Z��޷����P_
��RzG��\}�M��3�K��$q��HF�	���Qja�&�3;*�Q�4��+���-A	��1C	����x#v�,g�x\e�pꍶ���x�x�F19/���]��Ktz��ѩt��>�]���>�� S��P6Ao������-#? ˃$�A٠|x�Њ�9CO� i-�82�s�A�&�@�q$/0=oS(E�"�#�׵�7���J4(�W�a�-Fik�Gu��8T�+|�� ���:�j��9ؓ�m>6�܋W���~���	f��s��,ҷt��f� 1�-�m69%)�7|�݁L4em�^�Q��R�����������I���z�4�=�Vj6�x�~x���?/�CL'P{���?�j��A9Zm�ֈ�8_MQ��1JX�@Ἕ�,%�4�jv�\9�۷rl<R@�VY>�c���X�P���ǭ?�x,4:�.����i��5�>5���hcfDA`eϩ���������Pl����VkgM�6�H��E�aAUf����~�������G>o�}�O
0����[|0���Ñ���	<�z82�K@�dCz��̴~���묪��Hi�E�K6x�ߐ�uY�c��;)2��:��:䏱j��FX5(�=�b���_|�ƴ(
���qU&����3t�Jj^!T}���5�%��V�]���J���`2G������-j��J0��:�Bš$�,S3��s��}]b�O����� +�d�Z^s��\�%ۿ��P�:��d.��,C�})�������i��U3�r��j&��� q?�֕e��F�Q�1{��r���q����B�� �ͧc(&�u��$V�P�#��C#+nN�g ��3dֻ5z[`t���?P��7�]��$�Z׷�n�&q���*�P�I�D�S��6]��A�s*0�6�9�����h5���\C��8I3!#����ij��[�K3���{
�$�+HUÝ���1{�*�fn)��g�H�'�s������T!=M&�0�Q�C�5��ƚ`�����<f�/����Y_ة�3�{]�c���M��)vÎ19_AY�n"�~�2��-����X����4v���VӶ��\s��6�(Fs��Ϙ���!䲀{���(�D-|kBZL���rW���o#�4�����G�לА�dS���_j����:=�~�5�'���s)�g��9g��I,���rkD-�5�*[=\er��p���X���!��)��wC���j�sD���_�<�  ̗/�r�A�O��f>�3?7\�#{��_��I�]Ӝf~���> D��|���>���k2�K`�*S����@��MQ 6؀FTc?� mں�%���s�L�Ѯu�$�p�˟���v��=ȇ<���ˌ7�p�{
-��:�c1/��?��w��d#O(f~[��
b�a���w3�JMT�<5��z�(�'~�6�`om�둄Kًщp5]�^����%������V[�+	A�:�*�l�F5OD�M��dK��hN1l����*��7>dlЉ,���ҋ|��~��VYȩ�p�����a�S���rEp�g�ʌ���
��������V��N���"�{IU�=����l$ J�A�y	�!X1�zqM7����(���u�1K���lv2�X/?�ԕ�� �k�e�d:,�[�v��N��c^5�Fg�T���S�Q�n���m���y��:KRS<�t���"���~���	�a�x�0��7����uT��;�#rݽ���ium��������7T��b��S�Z��>��|4(]�sk;2���I�l?o�Y���20=��U���>e�t�Mb�%�[�yT�9��K��G��]�*��RRrY�Uܿ!1��RtB
�{�>p���9����[�fݹM�N��䲟��-Z��MY.F��G��H>�����z(� [C�����q@>�M�Q{'U�tL���a��-���U��� ��h�%���^-�_����
�����3V���������%D��>��S;,�A�ZG��~���X8�5��p(sc��|Ǜ֟��������,q(�q�Bh(��m{Q�7(���܋�Qup�=���j;���'���)�,���ߟ�������|+Ks��{��\�V��GQ�ٶ�&q�8{0�@+��SMO{�7������'��<����Mk�C�F�������ɚ(�J&��X���
�y�H��7�D�R�O�w�Mr֐d�L{ثwYW���������H�xd7e'�qHg>��Ό~Qo6�D��%B�۫wz�Ԁ���jY�VK�H�����ϋ�M��\��+̹�(�;�Y���j<��]��Q�8L�gd��	���t����4Oo� O�B�c��O�f�cr�}0��Ra�%�C�V�|�D(�t���d�ʴ#~ܩFLà<�׹�o5n�`�/K���z�&�ݛ�H�H^�ѳ
���P�p��yx�3g���侽(>F5�ѤFQLg�LD�F{��QH���2�$�G3�:ߘ���CZ�S��?�*�L؃Y�p��"E�Svz�ș�u%��<�8���O���`����g�'G�9O��_��W��1y�ypY�|�tE~4ollwPL�e��7�o�9T�s�"�vД+�ʛ8�*|I�D�~W��?#�N�6�i l^�a~`��\U"��#�NQ��$�x��s柷(MY�{3@����Mm�S9�����Ƿ���¡\93�'�������)���d4��I����N�{]3K]1��E�%.Pۘ������m������=bZ���
}�k�[*O�!�G��G2���v TT��y}�	��Ӵ 	1�кen���,U��!L��Ȫ���X�V�G���V��6B[*C�o��Ewv��[ر�%���^���h[aJ`8��Z�I|�= �4���j#DQ*�?A�6�����������z�0�@�9L�Ҕ+��pOĶ��b~�	3G�v�^h��C��ֱ�NN��/.X[�L�f����ˋ#��f�lYng��k�����t�`'�k]�i��j�Ls��QzG�f���):N�� �Z���S�,�iE+^Lt	Ya3�%k��#ւjű8(0��� P	,���3ɼ�9���U���H���A0�J3&&���� �����e���쳭U�*���4�J"�c�+�wI��4�D��s�P��y���J�e���qM��K	�6$;T��7�'�I�͡�f������"(��P�LL�mZp!���O��O��O�N�f�����H>�uRA5h��U�#��^�򾞛g��(J��'N/�;>���鈃���<�e:Itk3��ʚcB��X�5�Y�-��B�v�,/+������S�X��WKq�B�sa ص�x�3O�\ �A#Nu����[5���߇����!)['`�b�Y�DE+'��x����z��)�=�
��\�`��_*)�l5GҢ�{r��,��
� �ܜa�V��P�4�X	���ks>���2�}N�쿲m�����ڲ�|Y�W*8�L�I.��4!�W*����oz��$�E��*��{=d��,e|��4��*�պ�	^�-J|�~$�=���V$V�H�1�c��Wj�7��*-]��eo�9�.w,�����1 �Cմ�����/���5�ik��M����*��j|��^�kBXU^ݵ��U��E����=˚�˟��T�;|\�T��!������B�����~޾�t-�ҁ�r�����tD��y/����	���u��������jݽ��ۿ9��?K[u >0�K��(�� E4j�ɢ���` �0z�?�.S��~�o�W�;8�P�b}|��+������n܀��I�MU®��z�����"���MZ�����}S���q� b8�J��y�HzS�n�&��!/$2�Z4���8�>Mq٥N���@�b� |�w���/�Yς��I��`z��gJ+OE l�u�
�����Z{�v����a�TCʿ����#e߾B6Ҙ�3_��u�	���q��,�ݲ���œ=t�������M�jMMd'×����]��2~U�t;����G������B\H��k���55��Ƥz*��7ۛ{�ZA��-�o~r;��Sy�0��Y��)&}�<���Ǡ���狴T][���P{�DX�^��!��w	�f�$HC��M�����j>]ˤ���ԃQ{���og���
(Y�&ّ���sh���md`q���5R,�x�s�QOʑT����6^+0�8҂�Bg��/���-[AHJ��>�C�l3��8!�6�{�(�%�bG�І�jG*��`��z]�s�h��r�@)��XD���r��cs\�A�y1��� 4n��-������uh��6�A���)�|5Ou��H��kU���*#`(��\�xe/`xt"��
Z�ӝ;���c���Z�z`.O>�Rg��1�׵��me�䫪����/��"\X��n�l���������� ��5O]��l��#ES����>���z����g;���BV����	�)M�v�\-�N
�v�����<G����M�ܹ*vg��q[52�k�*(�����Նr�8;��87��'�a��*&�d'�Bw��-h\��Qx\F7�{B=�jgV�2�����}�s�(�B￸9�*�Bd��{����b%�����F㘨)����;y˶l�)���*��=mj�,�Q-�:������o�2���7ƣ��j;�d�U,�jS /<E>�����P��C�,6s�;�I����?�18�Ax҂w��5cO`-]�k�.��&�z'Y"`x�Lǆ?�/�8�Ľ뢝qLg�,Z~�]��X��ɯ�.V:��5���F�Tx�id��!~i�S��H�@�� sye���!z_�c-x�u�lP�O�����Z��	��t��gV�h⟞oA~ .��GL �l�ioM��y�9!�$��xT��kz�bʓ�2U�ظy����ю�c����Pρm����!�d�H8z���z#��@$z}X�QǡǇן��\(�)?���jqi��8W�'���HQ�j�^�0�i�)�~�`��g5�$(RM+'�Χꑯ�P��=�s�E�՜��4� �������Y���ʒσ�0��%#��IHC�l��x.�(�������s��aj�Ob�P��#Y����xr�9u��2�[�(���ECj-���!0	ƞ�-�pW�T!���sú��Np�3���O�ޱ��8i���t�%����cZd��gS?���P����j�*ڧc�D3�x�G%�)��hv(���.l�ب��ѕd�n��?��ȺC��|��Z!������-�0ջ�
ֺ3�0�.��b��sIL6���OG[�~��1w��z�����������;S��_��4��#]L����i���@g0��� X�Jt:�a���C�A�^3��!�1ٛa�f˺��9`XY���]��F@S	Y4:̕��_���@ܛ�vT���!j,�a���P9.�@�b�I~S����֠����Q2=�ell3f�$��؛�M3��c&e�:�}*���=�>a���sK���1V�Hx��j�UC���u��
���c��ol���%J��S�r;����Wy�ɤ���V��h��K�gCw���I塸���f����d��n���� �T[����	���<0C��F���t���TV��ݤȧ��!| K̅tԖ�sjOt�D�Z?���ʹ5
���]M���I\����w�+�6,l_	��$)���;�N���?Y��פ������`�!,���|c:.�u���Z��Ur�/29��4|Wn1�,S1�3HGT�=�wВ���.�xss�"%-�4�zḬt��-�F-����}�ph��T�{�T���7a ��k_M�Ҥc��p�(��ˮ;K�J��tķ�U�I����U+N���ѿ�B1�ϰ �K���1�܅b7������=���o]�h�=1w��g0�����q�G�O}�?��J���[�J����j�R�,�A���|2/������S.HCG:ҥ9���r�!m�0'Y��E$}_��&��p��k�"�Ӣ�\�ڏ5*�mPQv_⬗��#���D�0��X!Lo��h6����3�Z��Y�FO�AD����>JQ��W~�[¥�o�gl��6N˗WE�g[Ed�lsvx;vu�_Z��JLP���D
�h���5͜����k��&����Y�8>�ˬ�'�&+?O���ks�e�6,�^ ����+�T����tj�S�q�گ�w��j��Xu��r	�s�25�]é:��5���ذ�N�1�3�����zW]�+�O�>�'H4�5"�kR���bd'�o�J������6۟���j��?Ф�S0��:ʏ�Br3�c��2�,ը�ы>?�".0׺�pԭ0ޟ��7��)��ܲĎ��fi�J��@�\	��
o8'|�B�z����ِ�#����v�������h&�^'D[<o<���kt>#`j,�]n�Ə� �+\�=3���\��C��@��N�.yЍ`j�ο�;��R!���b��ki�J9�����
�Y���̵���~�:In^��j}�0���}YT���s6��J�	g����S'��E8^6J
>@Լ �{��ir���{�l��:��������Q�d�^�*��I��h��oU���I���_����V���/�:����W�޾�k��\~�>���u�X��^��T>��6R�!�O��6Ia2liP���ҳ���Ζ�mH��U8Ϫ�Ƿ<���?�֘9�ZT?�@�!�i0&��N�`ȝ�cT�O�RU۾�KΛ���9���Yp�1�}A���5/@8�]���E�e��^�p>[TR�6�X^Ň��+�7Ǫ�Zs$���j�;A+�?�P������8p��"�i�ۯ�nľ���B��Tꌥ�WN���GP�,�Ν�d!4�YE��H���.�8i��À?Dmxp�%}R+��xyX�f��}d��lx�CŁ� ^����x�63����Jm�*F�,��vn����(�-Z�e.��A��nĆ�EZb���P�,1�O�Q�f������׿;��qHw��&.��O�� h��zn
�uB�
~k��6Ѹ���V��)��xF���i�#�MFq�����OO
p���ބ����<EEW���ۭa��E��nm�<���NXW�r
�p�8��T�Πi���!j,�,�K���)�R�W�g��Dq���HN��sH�&:ۚ�����'OH�+�?�Ӻ���.�wΔ�b�5f�_��eB�f�;Nm�a:D���!2�M��R��v#�lRYu�υ�����f��°�y1���65f�(�1^=�@xz���d[���J	�5�F�e�ʔ`r|����\�҇�@n1Y������i�9*�@�;>����[@in%�H(�o��ULL\�a�I��pߨ.���0�uVª�>Ѽ�B�ً�qY���*��oD�0�QI_�
�ui�~�=�֑�hE&)t89�a�I�2.�~M[R<OZM<0�Y��*�1�����
v`�x"`Tp�av �^�ڦv3 M<��w�m�?���@�KF�[��c�t���)�Q������]&��E�u����u|{ܵo��~P6��+�1Y��s�����.��i��Y���QqN���򔶰T�������|F�
V~�媱��a?�CpȤ��Meq�y��Q��D��d�TJ �0w��M7�����q�Mp}��@�� �C��/�L��b��J)���L�w��t��^�z'-��A���xB_��o�Wv,)e�29�ٺLa�~2��6����x5�j�g�����M�.���z�-C�換[�Ν����3�;���G��V�_�N�f��>�I1i��[{�U�ӧ�v��A��T���u�;�E��U��l��RE?����-����f�}H�W�����-�q&��Z�*�T��$p�b����b+T�A(��������^�QXbc�r����히�ꛞ��\e�rhA�����&��K�k��2��*��'�O��G��{��(�D��9�ۃ�O|����O��V���lK�e��\Soʵ����"����-�����{��.�؆�K8@��{5O|���5�?�����T���2���#��6�Ϧ��T����F��]�b=W���`|�f���>��
���x���:�Eǩ�K�o�؞�S�(�����;����Mַ�6���N�g�u���|�y��ݬNzԉR*��� lYǙ�h.�
:��l�A4�պ�l��� X^�E�|$�I��+$�{��1N��A(v�r��ગ�H}Y����^UF�E��t�>(�3�8j����B�2bV%,`%P�F]�O����
v.������|�T��U;+���Z/��B���o ��Få��A�a7Y����:�{�VQ럭�� ����<^�Zܖ�V�y/��*V"t�?!���34�����uQ�����R�f}v��@ˢ)+5�=�ﯔi)�G#,Ro^k �Y��y-ݍ�QW> �tω�I�d	��ϽCʪLe>���y����$v��(�#6� �����=ȖZ��|��6�{�mA:'a�r_�li*~����2]�^6CJu��U�س����d��sNѣ���IaaY�W.�D�Hd�ئ����14��іl>I�s�,Q1�@���UK�'���"�p��1jR��2y�X7O�w��޺84ɼ��}��N���ʭ�vcE��8�ݛ��>���r�yRr��3���L,�<|KTI�U��5����z��L��"��)����s�Pt��0�
���/
S\S����5���"S�����_�����@����#g���)��3O���r�'���|/_���1TF����TO���~'�Ij'�p�ȟ��K�qH$�4�f��ͮ�Ó_�fX�E+���)��i�r�<������Y �%�;��(�'��7f���0,ÿ"3kj�����F����"��0��;��P�O�ǑM����a�m ����
��D�R�w�-�o�e4�r1R�x.L�����-��1� �ʜ6�@�����}�'������cD֠Q=�4��Z&��@�싫Bn�˾h.8
P���>5h�
��&�������9����\&	)�+L�����EzS�Ϟ6�G��g�}$C%�M�	T����f�D�MC��|�Dl��1�u�|�e�T�|�@�=*������듞	�ƍ��� q��b�L��!�9a��#&0���Y�D\)����b.�6.k72I���TE�b`˷��怛.�Y�Z���|dR,)ą ��A&��E�ޑ�&n;�Z-���8A�4��^;r���2�mD0���
ooA���m<p_���ue���0�.��܀�t���c{a[D�O�MԓNH	�Y�3)d��6Z��g6����s��svPz�$�,���a�IM*��z)���R]�c�3��|q!�Yk�k����6�=b&Gq��:F)�TRJ�ܵ��2e,(7@	��}���R0{OQ喼�Yk/�M��^��ԔK{߉w^�]�Kh
��G��� �O�:n�0-�����~q1L ;S�e�8�d�G"�� =����a�qn��V�u',hh�D��߼?�������N|� ��Xf/��P��҄v|�~����d_B	N9��V��x�~|��o^�`�}&0��4 b@�����v��HG�~�@�s$6��|�g��E!w@�>���"�}�~<B�l$�����z���s�9�&2N�͹�-�
mԔ�/{��Z4J�ʲ��Ѭ�xs��0��� E�	9c��3��行F���tɈ6�/Ш1Ͱ��SW��������X����EC7�x��B\2�d*W��������l����H @�qe�m�²JQ-�5� Iz�������2}��lH2��{w)
&�gyn�h���c�02z!�W�f�q�(�;VI��cE\Yx����!{#�#6m�9����O�k�@�x���d�a�g��.�ڙT���(M��Y���
Sb_&E���	��
oy�sv�Q�]� E�hk�9�����i�Ɩ8�I0;oem�m�d��9�z��܏"���K��^6+���W%6��А^�`3����I�A��>T�P��h3Jw�-.^ܠa�sh�Wx]ܦŉ	��ߤ�2�����T�6�0�����'�)�a�Z��|H��Z��+ڵ�lP�v1f�䁻�r2~��=e`Gֵ����&/����h#/�)+-�N����J�Ež2�����ZG��Gg{���M#��Α���l rZ�������6�Y���p�ބ����c�35�̷���鄀ն.7�`*[T��i�s�u��n����yT����*X�Q������ZD�O�`D#cJ�N!��V�ų'	�sƋl1 o�x�E)K�C~U��qi
&&q��O(�$���50� 'E�����mG�V�7@!p���LIr)���s˻������.�t�{.��]OQq�S�^˨ȹ/}���w�?r��t��Nm��+����!� j�IL&����"��4�D|Z�4���d�m�R���B0�k�������T�9t�թ�tO�N��u��xG���T_��%����X��\Fnдܵxy34��NR@uU`�շ�=eUo��W�o�%ݚw��>����"���E@��aQX�V;"B��[�'�$n���e:��9D��Ŗ..s�N+�L����
gO�am�	���4:#�~j7�K}����?��!���[��*�͙��.���^}� �k��MR�Iԗϩ�M6��;&!�Y��w����)�X��f�OgJ	��\�WaN���8��K�yQ���BVbz� �p��{(����?B1�7�-����k���-mGE�n�d5�uN�D����� ,5ǈJ�'IBi�E�)GOȇ��u�Ʋ�M$��O��R��$P�5��Pi5%m�/���1e���|Fh����^`�u��з��)�<�m�s��UY�.y�C(ًmZ�Êe��A�N>AF���ij��R^폑m,�������xg 
PH��������sJ�,jW�NB����i��=E	�h2[6�S�Ը*��y�?�<�����#v��g�o8o�8�W�%>5.��>[_ڭ��y��YI�ϒBE2��!	z���N�f8nG.1$�$f��[�In�1��r�2��G{y2��՜�������V��*��=�i��f�9<}��S�U�(����I�W@��m]TڌP"b�����;�;Vv�j�����r�k$	���C�d/�٣.�	���Ҳ�& 2�C��_��^����j�*�[�Z��y)֐n��A�ĵ48�ߨ���Jw�Bh�"MΤ5r\�[�+d��+��~���?��II�/m��K���!���n�h���ҵW�kFf�PV���_]�@��:M�і*Ms,I1̤J��9!,;?������ϊm��V�z-w��-A���Č���!H�Ḇ_��2mw(l�����:�ƙ(����k��M*����Y�����Bz�<N��?kVbuu�}c�`3��o;���bh]K��~� "<�G�Q'��e��u�57�G�e𓜹�59c����`f��J����E2���ң�sS�2�i�Z�����)`:K��N2��������a�]O��"&��5�r��5#������l��ܿ�(�>oг��O��LQ�V7����$����,��UD�#��Yb���y��S����u4"�p�0t�(������%2���!-!�)�����Ǝj�-�F���'�S��ק�X"�*����~o����+]�d� ��>j�=�zֱD�_h�܅�I�|�tw�q[m1DK?�L���`�ׇ:<���j��M�E,�P�N���\��5{,Y;�.`�X�3�0�x&z�}����N���/�x��.���.���Iw��_
����q(�������6lvk����+ۄV��^%�Vs��
;�����A���0��/�@=��?����9.W����Ր���9� ����F�1�bb@A���țߑ��j�@H��o�ٶh�dEg�FyW�}�
Bq4ʩ�P1�jͣ���>�\S�yj��B�^0�(w+'B�Q)JΏ+T$oN��bo,~���kđ.lƃ���Y&yǨ�n
�z٤U���@<��Z=��r E����J��GIK$C($��W�d�K�>	7��g\��]g����� �u�-���%Cp�M���W(��-6��s��qm��/������@��t���/5��J���W��MI�M�fi�u�f%q!�	07�p�]�b�T��.�EN?>�.��+�_�����^����=��(4|>H��e��_��xڨ�{��k�[�-��0��~l��_�͘�	�?�R�N�J)�!�QI@f|b�O[-%r�<79�b$��-Q �,����i r��(��GwKu�-�@��ݕ��&�+�`��r�]Șt�$x�ǊSô��L`�GRj(�4�b���/>_�s0^t;��i�����iO�IKq x��0B/�{��M��A!2���s045b\�s��Ⱉ��5'�"�i���*�	��$��Ppj���^����[�<Ӣ�u�i߫��k�� ��!���r�f���J��iP� �}��9�����ZVoj�@� ����`�h�"�ˣ���t.�9(��B�p���Ϊ���E�+yl��T����gg#�(&�xe��IG'Au�@K��r�<�٧r�e
U��>�%����]�}���B�:[������� �Y8�9�Os��(V�� ����}�H@C�Wx�3N5�NiƠz?�7m>���47Q��cfD����VM�� "8�#�eNU��G�a��n7-țZ�`��o���+6���|��[�C��w^:��u�Z�a���)<}3ذ-\���ֹi�_'?��2��n���G��b�D��Q[�Rނ�:S;�x^�sK�ƥcޒ���c�x��l�VP�e�@3��~����w��������N��_����Ҏ,�_Vavz
83&����ED;�K�}�C�lYb;���7W�+GF��8�m1�#wTk�
���u����O�RyM�܍J+�ǆ0�6���s�ΐ	��"�Jŵ�˺�@b��"���:�)�Uq  ���/�aL�l��g��U��z�j=������A��Ex�����t,����Y8SO�K��d菱Pzra$��k�	���Z�OǃY	l��[���������L��ҷX�x�=w�޲�H��q9ß���F�?����OƵ�6���?�z��p���Lƴ�)2��ً��fh�P4�g����>��v��'��72%Ҭ(��v1O^��1��Խy�׋��,7]�k*,�����3�Vl�0`���%�h��J�NX�n���?�k�=��PӤQ�c�r^�ZTtAx���#�5��>�(�������~���J3�g��oM���=��/�2R����F��=�� (2�eJ�T���#Jƕ��밵
��ϱ�>|�L�7i�l*��S���_���M��ܟ����(RVzo���`���u]��}n�SI)�^3ђ��0��q��>���ιć�?:�u�r�����|�����#l-w�~��Bه��ɟsaa�����S�V�y��`��d���c���A�	w@�����(C�����;a*T�2��؇K���1o��=m���C�V*5��)��A�]��a�\�����^#9�L����3xy�\�_l{ŧF_Fo85�6�q\�Í>)IE�Հ���eu^&Q^].짯���r� ��?�:����6��P  �rkT�Na�Ei���f󰫣e��
��rb V(�X�L�<�����k���0���<y� ឱ�K1E�v���:����⁙��T']���{�f y���̛�1;����*���D���$��=ЬTX��U{��ZN��b����$���T�4;���1:�y)#��$X�{����KH�0�3F��p��*�����x.� ���G�d�@��Pi@�[��5����B��/�&�g�Z��|��L̯�;��JX���$G���ZH�NHNQ�~[P(vs�Ȋ�'�c`�r�������=�Je�\��x.�Wb�Ą鎏�u�dn�h^u��<��_�k�$�c�$ �U�@Kq��̽T�2���pJ��qS�\��9�ׄ?�
�d5t*!6���-���z	��Jي� yF�( �[����\���t�N�S�E��{E�M��%O�b�����i�W̉�/������4���w0�g1i�>v���y� d���3�O�U�?*ܿG�m��!�*93@��Z��@#�Ș�M��jg�#
�mz��j�C��T��q�+�
�O����@m�=8�#�/�.�\:�E�<�*RN��^����k�L��g����?�ZQnv-'30�Ok��g�7@k�T�Z��妽PK�O4We�U`����K�UJҒk:��D�4�^�ԁr��|%����xJ��5T^TB>����P�,�v�ݞ=��B�����z�aU��E��w � <��#�^ ��ɦ�'���*C���?�c����4�}�t�1��"c�B�Ϝ�Om��3X�c��!'}8/�1(<�.-�Fe^��K�;`��r�:�S�-"t� 3�"B��>�hyT��
�e�)�f�d�q��r�u���"9y4(�]�Z�-B�nh�;��%��t��D �{F*@3���8k�G+/o�O}4�i)1�݁��܊�����`b�T�u�E�\t|�Π����L�^g�;�J�.��|�Ac�yXԤ5t�m���~�� P3�D��M�^PnĊ�K.ZE-s7�(lޛ��t����c�q���b)ͮ�w$[I6�yj�}>"O�+M�9g<�Hܧ�D���Y�.VՃ�y&�i'%'�9�MTHv������ �?����u	�KZzv=0�{g	�Y�k����a4P8�a�Y���o8g{����iV�n-�(�f���8��ٰs��o��hwZ�
��kAj�ux�0���<�&���i �.lĈ����i!0e[X���_������B��.�#�0��G�iu�aY��igP��QoR(�y�;�TT�)xp����IPL#����x;С�Y@A �ړ��c��e@��ܥ�-�s��3�##'��RQAo��� �=�2���G"y�eՁgJ��o��ŏ��c����U3�b3�m�]���G#	�Dq%�jZ�����	�I�FA&��%�M�������<$�x�����oO� H�W�Q)/�*5<(�T���s������}�sp���_t`�?4_GqT{t�&5	�G�ת�3n�_�@���W�s���h|?�F=�#|�k]�&��'�|P�s�(ϹЀPg�+e^~����n�=`��9q��%���?�O��]ia�^Q�<���⫳
2N�$�K7a��oJH+}t��ܟ�M>$=��}(���P�;��z�z�5G��� �!(<��pc�Ԟ ��}�5�jv�qk\b?�$W�i.M1��x����̂5��o�sh0��ʨ��#�x�؂��?A�TLɋQ�&�M�5G^�@�_�%π��%���%s��؃���)F�a�9�[2as�m<ӗ���e���sڜ�i��V�d�ax� e.���"��".OfO8�?�b��&{��F�~���mk�[��I_wƾ���f��E����b=�*�&N_w����'��M�"���;�Z)���ȆqD�D7ۉ��.��2w�y��ą�*>m�7+�X(�|�mٶ�=<���2G�"nXK�G@xOڑ����a�Kx�*C~�Xs#�h��$�ծ��c���d�����8��7�=�Vҡ���B