��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:�Q�z�n2�H�U��θ$ÊaU��mZ�^	��H��3��y6�B�r޿�������sJ�O9��j�{��J͕�l�q�"�dJc�e֮V�)`��N?J���5�8�����+�Ml��(L��nm��ۧV�;����uѦ/8�:��LD��� s��P����}��lC�;�����"O�O���nXu��X���V;H@�	,/��	Xs_L�86GvT$�cW�	�.#�O_��NѨԉ�;�D��%��P�+�������c�Y*�����`e/�\I��u�zр����f-/�>+���� ��OL��92���ٞ2r�y��oe��8W�+U�,���l x�z�
9y77M���"�bި�W
�*������m��Ak{�Q����h� Xpai@k��V/u+Us����ܵ��h.ٲx �S�)w��di�e��I��U�ʰ��D���`T�f��t�|L[-A��-��בRG`w�@bѫ��!j�ͦ�`����>�M��9����A�<)����S]��+Yn0�=��I�$��>�:z���j���9�i�o���p6�/�Y��'���2�L�A��O���:�}6y�%iwq�T�F�R[k�X��>Z&5T.��Tu���jܾ�IOS�4B�W��.��PhN��nl� 7�	��^�����DsA�ƉX���q	����}�7�Z+ᚲxhjK{Q�������)�;���W`�������f�|jd�1�[A�����O�e�8�^��a�X��R�2e����*y��
ٚ��P�;
�͕�ז���D�V^Y�\��4��ձ>�QlP�?�K���}�ʊ
~��[ur�Nh
� 6���G��|��~��d����b19�Ȩ�.�~�v|&(��LZᦆ��Z����:c�{�tm���n��X���ܿ^2�J��R(���m��<�S���vIb�R�E+�z����>��ubY����'Ig�0-r�2){�PB�~"Ѷ/ӹo�K2�N��Z �����2�!}bl2܌���O!���kjm,|׵��]����Z~�,�rt�&^��F�Fy��xg����f��C6�u&���yN�]P)wG����Ꮻ��g�e����@�4͸]w��E�eEBs�N��u)5U	�Eܷ��n\[ {�D�NJ�D�=�!�&����Z�m�`Ȯ|���?��yr���%g����E�Nf]�Մ`D�	B�|���Xގc�5�uOS����T�����D�}9�/dV"ê�#��}�dC��W��׼��y������VH��XJ�do��z���s���nBU���gA�*5-xl�ز�m�5-�q���L���ؼ|�M2�l�����?��S@�Q��2���.e�L�L['o�Z+h�*a1[{ǨZ�������@�2���t�
��Rf��s�B~*����w��%痷gˇ�i�:��/���ǿ�/*�D��6J�̢ކAj�:��>(i�	C�B�����y��x,1���Hz��;s��aLˆ���DO��ƭ홏�P�n��}]m��00˂8mA�WXN�X�©������sP������Q9��r�[����}10f,I��n����_i\����+=P9�|����BM������V�Ƚ����l�}�&���w>���Mn!KJ��(�M���3V�:!-e"�Խ�Y�i�H��27�&�\�2���й��N�O_�(y�%��~�P:��XMZ:��c�*�K=��â���7?s�3�9�m��g��34��kV�z<�&�Wr�.px(ʲz�eSb&����K��#79=��7�� ����`1�� �a����VC`�|[ň�Vi��N�;,�D���o
�Wg�#�8X���		��4�.,T�b�Vw�`�=K�{�{|=�s\��z��A�@,�C Z~��X��jC��2K�d����
+4�O�MW@�Jr}��z��?���la�5jC,��k���b�G�ܣ�S(箻�q,J�+3m��A��ɶ�%o:��8$SIX�&��ײ����n��iC�zh��>�vs�}���t͏}�r<����d���2�)��#����g�|��T�C�xN� �b�3�pD���<L6%ь5:��=��L�"(V��<;M����T'�m�y2i���x�c��^S�A��y�D[c���G\��Ź����m2������c��M��G����*��\j7J�؟��E\�馿���~��l���K�_��	�����UR�jyD���yƦ��ֶ�n����C���6<�
�.�n�}�BĤ}"A�:�2����2QZ��Q�|�n���h�XC}:�jQ(��
ń�ңU]e�)���ai�Ak�������*@{�ebk���"��А�q�&��+�t�Y��٭�V;8Q�:��J�)#��L�E
��tx)� c�ۍJ4��-A�O	Y'Z�{<�Uт���\u+M=�S�[q�9���3��@i'	N���l����&�&I�b��-x�c����S�?�<��b'�YC��%K�,��61ѲٙjX�\؈��!������,�%�񲑰�\FS��9�|����,�d#�~�/��Ff�R�ڙ���!w���2F�������3#���K�!�d�,ڶ�F��<���t7�^��7�u��W{� ��yj�v/��*{!��H`�5�%l{- jf�}�^�o���7�8�1����e�8��ʖD���l�'��Z���P�X�m}V��>�%���Y�lunz�=��o ^�
`)TPv ?E�ud�Z�ބU>n�6�SU_���g�aB'��?�ν��O�u�Ew��?,Mh��%�2��wŜM��pc0��Own.V�J"� b�mb����M�T�h���f��.�K���x�0�r�hc�D[?��+v��Ț�Ջ�&n�,�j�v��8$��<��V��L�Y���|�`��s����>�p��r9���n�:ۅ�4]��&e�K{��.�{��ۖ26֨`W��iN�o�Ϩ��@�x�z��'�4V�=2�_��'��&�]�,��Sӯ$����^mp�&�g旃	�����H��TxF�q'J	���I�����aQGt>�~*k/j6Q���Q��X]B��Q�lh���}����]�0��B�������@����M+�/��/��ta����h�MN_-�c>������	Gi�7��0V�`nF� ���#�0�O��I	�@��C���AN��O)%�^�mO]+T��#HV�FE�U��bƵ����ꜝ�i�X�4� v�3��ٴ�[�D�1���ܐ'F@oǛ�=�]��;��7,��\�,@m|B�@S�t��(�R����~��5��bCO��i��v4$JqQ�c��	��l��7{�k��~�_���7}�� ��=�BS�ҧ���{!O�o_�#�yG��m�k�ȋ,ֈ5䛁ɏ&��*
����=�4�`k^��CQܯ0x,��	�|W�4�G̍�yu\�#�~�p�U�����d~l��'�ܲ9�$,�i�f��к�*��b�[k[�ya�:���<��w3f.dǿ�%>V2�*�y�'�H�
]C�c_sNl���gFU܃�|(����LQ��m�'�y9Va��#7�v��p݁�*�ty%z7q�a��q�����G1P��b:��qBy�@��E�у��ʊ�ٽC��3^$�w;	@�?vpr����k���<��Qĥ�<}G��Cÿp�Y��i2ãy��M�v_5�:R'zY���AUsC�c���$���B)��g�y�ߛ�M� �F����Q�侬3����b�F�	����K�n�d7�٩�:le����9�q�
Ya/��8���J�\(e4l�s�DK��8�'�ɀP,~��B3Ӧ����96��|��]�$ǌ0 ���c�^>��
������o�\��@����\$8�T-��H 	tB��q�iT�����3�Y}����>�9��o�ηN��I}[[�/7�̝�
'�M�C̉F������x�5wH$0��/O�lNi`��Df"p�a��´A8��v�"Y�>5�T�J����}\�҆طk�g�@�4�Ȧ��jȰ@z�>�r��=^޺I��\���ē)x�%n�c&��=��y�m��f2`��H;��gZXaPmW��l"1[ !��J����:���z�I���fL��d7��D$'�	�a�E�� _�tZ%Fm#�e��mq�@Zp�!<%<���s�=>U����2[�L��r!�d�A�}�Gq��M��+@a�r8M��!�;҂WU~��FJkG'l��'-���h#a
�t/ˉ�"<��=�G�6���a��S�ך���ʼ�7�]e��߉#��r1�Hd��&�ן5�q�����C:6�
YQ	�Cg�_�_{Y�m3F����Э���a�-��:�����p��/i�ջ彈K�lEW ]�sa���_G�xP|z�9ȸ�8o�1��\��ώe�c<M�[��>R�BWp2��s�!�����s���b5oga�*�N��bj�rn|Q2
��ϻKzgAѺ�~g�Ƭq��p+���I���������S���Ɖ������-'�ĕ��>�����:�����4=	��h�>1��P24P��Aϙ����\�$g,��|�ॾ�1�^�Gxx\w�sH��]��j���m+ߥ���F�2�(��]�|���rGOK;�401��{�"�v���c~�&�;w9/|a�����Y���ޔR"��Z$�Fj���)d_�N�6�0��mNZ���ؽc��FZ`j�Z��D���9c���U���
�N��[4ZeyX�d�w����Z#��7��P{��"қ��f�8�>����|�
�Zh~|��W]��@�4�a<׋�.Q&�*>a	�W��3f���9o�«5'��Z����Hn�e�ǧV�\�*/qx���P궝��k����
��x�����c����&�O �w���Ћ;���HI����0��]�L!�{�C�����bP��ECj�xp[q����7Ve�Ct��T����齹	�=B}���rG�����e���Ҏ��+����4l�<ƞP1�ZӀ�:����l[	��?r�* �Q��:�+�_O��oO)⑬ab����.GHY)3��R�1�|e�dQ2�M��̋+_����sK>��v�UAg,���,2���+(��Z+���?&�=j]\.j�$H2�_�Y1�S��g�:ϐ�c�S��r/	���7�B���j��{}�ۜ�� �V���v���� ��� iO":}}�F�UcpG4~P�'0$��J)��0c~���uAS�HG��Si�·���C,ސÀכ�ڡ8t}Y�D���d�C��	1w�N�N|ʹ����/��K^a6v�#H�۩9�]�;�%\�'�˾�;z��t=��.��<��Z���R�-v���,�5�'����G�� �m��gǰ���9Vi�ذB��4ӡ�g��<����Z�'�
H�Pu!O��.�"����6�C�g��&v��:�}��L��.4-�P8x �.ѝV�C� �\覨���C[�Gi
U��,09�+xu 1��З??�<�]���В��EAd��G<�s�_�+�������<�Ow���go��lz�ĸv0��k�" j�k��E(�2��5<�	�%c��&���A�zq���%+%�bJ:f�6���F�X� P���%���t��_�to��7�T�;;�v���|d6�}87��ޱ�t�@�`�$iX����k��G�7���[����w�NQe�l(�:1N�ߥ���Dwlm�<,��G��6����R��q#�U�VIw/T��L�c���W�	�>�S��x�������*��GRGJ���3�������;�s]�7����� cR5��,9].�O���{+\�#}O��ɷ�þ�����]�@��u2M99�˭C/�V)�ҙ� ���9f�p��0?�՝@D�����>��\* 7��DO���lI��\B��	�y���=����g0��(Ң]���q�����o�S
5H�Xp������K�\��JE�z��� K���o;�+�|eXz�x���A�@Y�=��"Y�k�S�V���,/�⢋��i�a{���S�W5���̃:�`Ω
�Y�^��jeJim��/�����u/���$f��9&aOx����j��v�L?~=�TP�@��)���\�_�sř�*�����Aq=]H�BBD�yn�P�~�Jە����7ܰ`3�����{~�gnJl�-�Y rf:ex�,�Ǧ3)N���c	����ú��A. ���$�:�t�����O%�C�Tu�,-M�,��ߗ͈��tA\ө�~K�U�ˁI��vZ�߿�q�D��)��-΀�LL'7�ֲ��5���h�����D1RNZ��UsK�qd��t�"F�E�c�L�M>-��s�x�(��Rʭ ō��a�10��\���;1r:/ĠI2oӈ;��"�B�]���"4����j5N����t����ԅ�tș�(��v[����h�"���{/��]���e���a�Y�{�����E�|l��C[9�Q�kۨ���y� ��s��4�2�೸�
�~�	R�ϋ=�Yǰ�-�A�R��������S��h��b��t�"�s'2kF4 �SZ����w��}v<�p���_��
q�.�,�%Cz��0��_A��� ő�!�WgCN�p-��dCg���
N{���y�I|@�$JIiu�?d�<MD�z�1� � J��~����#���Z��L�5>�*�ƫ��ۨ�O�d��,Ձ��|s33�/d����!I �?�0�����uO�-�麉[�ؘ~P�
���M��C��^�!gb�*l]�C0E뵘�C��:��U�*Lq���<	�p�;��]QL��8��^�'��	�>�S���b�U�7�ʍ|�b�U��H�����_��}`vI߶����k��:���}��d�shq�������\�������2>W�y��ɮ>��t�Y��B��<�
�1ui�*�f��.�\/r��.��F��]
��{���O�;([��.����y��w�y5��>~�`?d�Y���dJ�q����x�ظ����N�ଢyO�� ��P���J�c��!���q9|{�=�k�%�?��6�Tɿ�Qr������V&w��8�9;DR�Kx>��i	
^�a��{Y1h��n۱�;�oD���#�<��ey�K�]D���h�I��ѕ���*�Wg^�'�)])eդ2M�t��:����gL�q��L;�g�N͒W�R��UT�l�_���:���.x����b�|9��
�VHG+��n׿�Sy����l�k+�*��B��^G7�E{�wg{h�5�ߔ��iY�e��$�,Ǆ�0d��K�K�C:� (U@��.��n� ��O�Д^�Ӎ��
Ed�������:�ֹ��ñve�����3��H����۹ѩG�^9�s�Э�W�����o���r�pAǩ��#���G���M��5#ׁ��An�-����A��<��݇�9Ԃ�8%����;�Y@J܃��}2"�����쮆�g�݃*
����:|��y�0���6���Ƹ�\��H�DD�j�����>�є��u�#��?��'SQS*�-s����&g�||�z�;���~v���&<���"G)�a�w�jfs��2>/�,Y�vn�`11P�N��l�}�:��Wܨ��}�s�?����hL J��r�O�Zr������,%�/�Uz~� �j�e`��Z#1@�X#\R�-���>@T�^��X��*}��S����#%���\ �=n��Ӵq�}ϟf���莌05��$������͚�r��"�s�6XG���� �驖�����es3�'���4��T�0y�$[X��t��;�:�"4��A莐�c�rcgx�6d�����CT��n��
���2פ-�X��`� S�$*�0[�L'$�����*U�̥�K�Pb�÷5_#��	�]��/s��Q�uy5u	����
��}384�h�N�
I6�5��BU���3K;��J�Ϥ�=�s�ч��#�s�!B��Ӿ�/�J.��s�&k��u�I��Ef՝�ϧf�"���wad�~��]-xv�n$���%y��o�9�.�TVY�fX��lW��N�A���H�4c��kb��8��		j& �z�E�@���~
Lk��,��D�����
�ߞ"���u{�ꑅM��9T�+�>03 d2!��5{�+��2�̮qʟ�a1<�O��?`6@"�2�K[3�F�o���G�N,�9�h��\��$Æ�!�G�8��f���#8���.i7��́TP���+m�+ph���h2:�DJ�qa�&$�E���11	�f�E��,�l��k�:,�d��T�r{Y�^�!�%vD X[��ٽ��� =��
�)����V�����b����� ?��8#>���۟�z��}/:m�Փ�j}$��4\EB�:a�Z%Dc&�.�|i��z�Su/d�IFw�b��q����߽a��O��] ���Ɓ�L@�]�ن�������p@b)�d�v�Թ�@��F�fp5� �$,�w �Y������q�^E�H�" �U�UGU󻢇O�����)E�/�&l��o�����>/�Cdl�H�%��)o��rl|��\��KڗDݮ
E����כ%e��15;����Me�tǥ!�ĺVz��9����2��r[�S�6�"�J?�XO���
6L��v�@��B`����%|��F	j�����J�yM��<A��F���$�էC���!�:�������Ք��&�s����p?��/~<�^�`�]�ҦloBw�l��mef0��4F.HK߯���Y@�3X�w��E���kg�8�0x����hF���>�~d���h���)���\�M����l�!ƽK�m,wCCV�Me3`��#%�%~��4���uٌ-j)��4`1�ђh�����!��s�b���>m~�R,3O!�\J��J�E$5'ߩ�߷,�X��[ȶM؍�,/��AԱ'�V��S�S�]����VYL1#��1OGԊ�pq(D;�g�7X3![���5ϳ6�tN�9�۟�y�JhK��[ñ�0��#�e���>M�#%�i1;�[ClcӽM�m>`��s�f���؏��5�P������xHu�i�w��`�yE7��	����P�q�'ѵn��6�(��/�@�X���A����
��R#�9�(���r4��U���l|�����ˋ�>��/_��\�r3����Z������/w'��Z�@ �,-�Y�";�R�0�)�����e͒MLU<�JNPN�Ə{m	�0�]az�Kn�����5�Ua����Ф�:�-��M�x��Oa�BNҝ
�i���A:���	�S ��YM�~+����V��jh��S�->f+s<[Ҕ�S�oXzD��(�hG.V
�0��"��8�p�}!�V'_ǃuI��R�:������n��b���u<������۬�pu�?Fzm�Y�@ɰ8���Js��2p�B���i,�j�헂@�r�;�;E�B�F����[������[C���#g��_݃��H�@:O^�"��`���;���u�6gԥ�Y�e�5T����*��|���D�������S	������������D��]���}�+ORPD��G~�Q-�^Ԭ|��zW��d��?췟��G�Y��xf���Ȧs�.)��+z��)��2@�x��/~%Q�#�G��H�Nw��V+�9�����)'i��yjk�{��7�ا�G��@**
2騤=�!:�Nj5�1�=Xs'-��bNx/,�~��
��q��;;�7Kq�Sy--.A2��GJ���������@��ý���!X������R��:i����=�i�t48�0�:e����t��{-~,��@SX�eQ�ċ���6y�~�(��?�\ra�]����F���2{n���oV:�9t��
��F-�  �,B�4e�)�������!^� ��Ó��<d�F:��7�'Z1������De N���
j�朕m���M�݂K�u�%T�8`��$vY��������.1y���&�ņm����6�ם��S�>3�	�2e��X�FЌ�ÿ����j��a�A�e�Ѕ����c(���{Dk�־�Z3C�$�ߙh��MU�W�m|B�*�`�RfV�av�$d',0��j��U~<( W�}�s���:O�&����Ȥ�ly˪���3��6P~s��7z��~z��9���ٖ���[�_b�$��P�K�ا-�T�6�4<���}�j>]=��(��Gִ���r�U��h�2�	����ٯ�×따�(T5���I������j�w��3��Λ��؄�8��X��w��]����>�%��J����~�RC�E�W���zނ�0��Ŕ0��pO00P��s�K@����@���ݸ5�7����|h�=.�%�O�Í0���Ðr�i,�sǅq�S41��_�^�_�s�*a��I-k~���1�T|O�
�%���+N����ٚ�LS�Y��N"���m}:�$u?�OP��/䣡$����gU� ժ����	 �i��b�<����� �C���� M���J���*['E�Â�*�E��ǿ'l���3�q�?R��'`/�(�Qcu3��}��G�=/}�[?Q!�@Z<��\y1��uL����-�˹�ӣzA�t����ꆚ;AjKL�Dp�-����2�\7?�sU'�_X{�c���/r�(��_�+q¦r�}K4-]��A�_҄�	�����缱��hw�#{Ԍ��A�����k<��	��X;�YA�r�hC$I�b���E[4�5<�%�@�_m��v�Ge�?������Z�~
�tQ_߭�n|`��2/2Ԫ7�
��N��yl�N��19���٤��+&�?!~01B����o������p�#�dqxO�F�n ߑ�����I�S��\Cm7B���1�l�N۝nu�Y��l4&����cβ��l\���5�Н$���#����ȏ,��N��i9 n�mVc�T�"�ekC��H,�#��4In�1C!ߺ��{�ニ��y���+?颞�l5�/��1���h�e�#�_U�9�7�*��!�A7��*�Sq� ��u��"T���}2�\Oًcy���K]��磍���Y�����9�(n����������ξu&T^��΅�:%�����ހ�,�a%�	L4u�Bŝ�)��rȰ�u����`w�>۞���|�����I���?����
�`+��l�1�|�s��d�#�c��?F'T�H�=���,,gZ���B=�ԅ��p/�׿>��h�Uj]�б�:����v��N
.[��2v�-��1�JLg*Tx�|z�� \��<��"��չ�\�>�)��� �O_v��o���]&=�x���܌� X�,�6��I�'�������Ek�����f��U��C�]�a��������T��?%
wJ���uxv�C�|/�:a[��WK�(���$�NV�Y�Z�Lt8a���S)��X�!G�gy�" ��� 	�O&ҳ���f���!��c`��k��ٽJ<���%\*�߅q�ZL�+g�|���2ڼ6���y.1գ�����(�R`C���1�u�����u���9���m����Z��X�/�	ȣ/f� U���x@E'i�M�L��oע��Oq�
��v�w~��!����r�j�zP�:z+tЬ�o�E���NQ;��dhr�w]F#qݫ�p���"bB�,��`d�MiF��m�o�N%���od��F���OB�5%.��;���7�%�ɒܪ_��o �삉m���
��G-�1S���z'��=�`�h#�����g��Z���_�tB~Wj��x�D�֦I��Ǽ�@v�l��J <х=��)	�d,E��$:z�$�B�R�dE�,�=@�e8V��+t���l�L�k���o���U_N͟���x�8F���fFy�ͯ��#�7��YC��b��j�k�~�)��0"Mc�sɂ���El�[��T%&�l��3B�i�N5KE���~8]�Ҕ����7)�1V^� .f}|�X��� I� ˁ�t��P3�4u���6��ey�k�+.YE���@<׵�$U��T��#�zE�-�G0�0����Q�U��̽:��7�� ��`N��F�=�'N�a$�5�8��&��hb��>4Հe�/S���K��݋�@��Ò�/�Z��gG��n[^�'�K�� ��!vȹ�*y��[8���M�'��]>k�]��v����n�u��.;���1���nj��	`�2����bQt���sLSSm�[>��I�[����-��V�i7�I;�\Ssi2�� �{�e>��bK\�f��%,Q��"�֗8x+)�cŀK���;��9M���/Ѣ N!}&���j�:��?%Z��%M(�4}����7��G��'��
J��R��#F60\�H �{
cM�~s��`�c������z�X[���$l�!�zHƕ�g&���(���j���kV�sL۶ÿ4N�&��$�=�? ~B�+�_�*M������9��PF;�М+��/�Y��&��	O��6�b �X�R�ld�&pͣ/d���;����8JZ�Z81	d�B-	��ʌH+Ȓ�	�g�֘���{��Ǔ�׻N�Ȯ��i���aI��V�W�������Jȥ��ҋ�	z�!�0��1/��NE�0o������aa�&�F{L:�>��;�A�.�5l����y%������S�8-�-���xTS���6{;�W�oօ�:l�f�j�fwL��;�1Qi:�h��Nd���Es
������7��Ac��F����>*�RN�5���}��v��)7��׿�]���n]��l*j�O�ղ ��+������pd� ��[ժ����`�n#g�׈�؁��c+R��ED��&�UN�EF�u��>�?{ �;B�X�(cY��!�^+��G�߳&����n���ŶN�� ��Pr�1:t�f!�d�ꧯ��>U�{/�Ţ&gAՓww�G�I;�RtԄ�:���a@eV7,M�Y��\�w�| 92Δ�&9��ݿ��V���ɺ[|��CR��Q��f��|I%J��=.�2��$y�ya���H���'��h5::�Fa�+�ֹ�z�Q�re����Z�L|���6��E�!x�hG�Rc�y����uȁ߂?e@�'D���²"��6�)tv�1DS"�ز.����1%�v�2����1��_=�A��d���H4r0�
\�,v��Ƨ����3[NU@�����y�t�	e<Ix��)m��
�V�S�O�\��Q���_�ǃop�̟ �솢���M�zgjs�p�2$Ŋ�lI>�>�­��y�Ű�]�s�/{?������Ԯ���y�U�j�ت�M��a��Tl����m�;0� B=�)�xRWJ.ր�g��n��V���ڗP����B�<q����u]�h���lT�����}lV�)Z����#ܥ���a�V:��Q�#>���q�r5ΡG|���kBD��J��f��h�_��u"�z�y؛�	�Թ�?��y1��!��E�{L/�}ۛZ��vAf��lv���w�A$��`��F�z,T������ziv���=;�|�-�^a�_�*e��T��E>b{�@��o�0<�#�{�1�0��tgj��\3I��u�s��	���aF�S%f1��Ku�Nf��A���Z}����s���9,�\
=$��M d��������#�o��n3���P��. :�L�.��4~М�sӮ5�Y'9{��V�'sH��Arv�i�)�����0�|Z�`B%9w�쾞�H_��ɮ�������@.G^-OMk�J��rK��l�Ԕ��0U�����A��B���f��R���\7n���п^T��S]���_�Q �@-�߹ԀQy��<����t��Y:E�s�砟����T�Ly߭SA����P>��Z�E{EU�e��q���P'T�}/�B�F�i]�m���#�ɮ��7ecks�4^�����P�	3��;�����|nP=׎N������xb*�.#&��eR��	�<wK �s�w�{�P1p�1����2F*��S�����٦����h�{�D�HYcә`�� 8���s<�"M�Bf�K���aaE��3�$�[�Ϛ�p��X�`�z�c�邍�z�~�f�]��n_ Pl:�� |]|�V�k��#M&4LBf���~P�6���\:�awaLB�
-�;SԲ��I��)B��4o�>8hVuba�L�o���_3ٰ牢ٺE���k!�P��
F���p�ۍ�;r�����v�C���& �Y���4Qw'j����H ��)'����*�x�s]�$� �.{�S��Jmn���!G�}-�
�M�\>nq���P�B�m���*uBU@�~�a{}e.�-�V��D"��\�T[���prp�6��"������N�T(���r�k6�-�$~�hp1^b��QZ�5;�'�=�d�P�XZC���*��Znj��_X��y�.*N���x�+5�!��9�e.cMr�qQ�,̯c���TR�{ɤ��S+P4z��Rs�`yb����"����'�k��� ��Ye\.t-��`PQ�jciO��[=��5�S���W��-�'�c����.l�t��/4m�b��;(�?��D�	$�~rQ_��Th��ѫV�_����4INK����'R8��'�.Q�D埓��A�à�=Y�4LBp2H�Mbg��ݜ�����z���@.g��A8j������uĴ��<�9c�f�E�yV*M~a!��@�MP�H�<y����>07[��rS���۷X�B�([���P��Na�z_6{��䆺0̿�|~�8DY���b}�#	�����.쎾띁+�\̂��aj�ጄ��Ċ�	�GoӪb���q�+21��w�g��Xt�dȹ_nӦ�C�a���̱n	�O@��8N�� !����m���SH��ڊ}�ɱ�/��,6�R9�%�O���֓��"Gc���C@����[�50����E@�n�ڜ�o���^��nH�����J��cU����%oϿIA��?����^��lIR�K��x|*_H~$z����GJ� e�5?��r Tw��3y$Ċ���P���g!F�Zq13�4F D{OV��nj(�1�.�W��J���Ga4�UF��5+la�8lU���Y��3��Ng���)]���i����v��y�&m4Yq����m��z��d���}�@Ȑ�D�K�q������l<�&H��>�[�L*]��)��I���q�Ճ�,���χ�+�L9�S�N�<`���^���ua�$���Em&�T���A�X!_<�W���"*
o�5>"�d�<�p��
�E� 뷚̥.�4ͷ�+��gk��,̣�'3üPV�>Krû��5�A~i�g�{����3.+��bC����T"'d���ꕈ�4�&�ۥ_��0�ĵmx����+�r6ǎE�h��O�����!R�ט�05 V<8��`o�ܮ\�P7�j�ݳPʊ��j� R�9�U�G�29�>�_
�?j���)�̗�+үr΅p=b,H6m$?!m���o��+�j�kX�D����@v��2y�K|�4yh�h����콡����i!�M:��_.�D�[���*x暎����ı�"PT;5��y�e"srs eJFֵaz�Q}��0!�p�w@7�.���<h�!z���|�fN�R%�v���*#f88�Iɧ�곳-����P)�"�"_~	1��;U;���=��":R�6˦
����E���˨���j@����O����� '�#�C�8��&ȧ`��f4bM�"���˾�s����G�S&?��곈�j���QVpL �B���S����!���o汫�I���'���O6�.����Q(����L�Ġʬ�g���(,bi6TdD���@�q��U��~:��=�@���z	�aN/�$\�oQ{�g��z�F'X��>}����� o�I�l-�o���5�UB�>=/��l�RDY���?�Y,7��\��B#�Z($�6S=�w�Xpr�_	�ǵNQ/$jnzKb)�r�B;�d&�����R�Y��æJ* �g�6��K��G����Ȟ�@�%�wSZ��;|�5Řj���:�ޓ���lz��s���2;�d;�������+��pz+ڭ���x�`1����c�/"������@�NV����#g��lW7�O1@�j^^2�7�,������g�_G�S�1����L����^�kLf��S�*�<Y��a�C���0�vl�es���W[=F|��"�a?��Z��1�0:��&
����<4�x	t!KIi�S�0�-jQ�MىX����'s��O�?.#��3����@p<�W��(:��W�q
W+�Xɪ��5�aM]Yp�ϼ��nC|�P�*�n(��:�>�H��������
ӏl�!��BE�zN�J��}�����w�E�7G����o���rj�ֲ�Oa�.q<��g&������|�g�
	�Se���g����!�`{�?��#OB��t�����l����E��V��i^����5!{��&�m���̷u��=��*IX���}Ur������(�PO�FB��s/�s�1*#5e��w���a�L��ɩ��ƘF�;z�(����-|{������z9��;5�V {:2�|��~��
�x��t����V��s0�0j��]CmK�1�G,k p,�:H��^��|I�XΤ�ϠC=�g=��	u��zDU���~~O�M@{����3��Y=ӴEUr�^f�(��K��v��ى7LYb"*/�}
�� H�uO�MHw���I�"�$Յ�V%Pl{���3�Y?��/��U��q/����J&�j��B��6f���SFpm4��F���E.��ǹ�xH�`�ݱ�����q՞��W)K�zx�>7ס��}�F�J���b����zI$@fW��(��EF��w�����,�1�Xpމ���V�G������j��{�ʯ�#���d�2�*��Z����|D���g�_Zc1i��hQ3lp�B���V~��Q$ƅ[�B���̆�E�H���sV����y_DZ?�h�!q��m�xK�Dc+��I���c���*�ox��r�	�vJqxH�Pt���zL��S+|�m&,���ۤ��h���t�^�aD?&z
|Н'�4�w.�J� n�@�c$�6'�!r�Br�V��|ń1蠜�U%��i-����u!�ܴ��3�k*�X/����j�g�
�\��]ZnW��8��X8�����4a"�pա~rz\�;���W(,����q�h~��<��Z~n�?��Õ��x��&6�{-�N��Q��y�M��MK��O��=�>�8�dO��@���*7%p7r*}a5u��ˁN�@>����$�[Ì��&馩��������]:N���j���ҁe������ea��P��5 吩`pYϹM8����,�hWڸ@������N��R0�7������`���_糀]��ݻy� BGN�����ٲ��kx�\����#(�_m! ��-cDkޒ�zY�~`b:}�	�~e��-�����o9��(�+�)����e'��?�j�vw	��v��"_�\ (X5_|��n"n�o6�r��VIA��I�����j�.�"��K�^䤃Iץ��)EBr����2x��&�vP+oDh���)��$�Wtd'�V׋�w���l��!���Wc:>���NZ�����E7�P&�)@��B��w�Y��E0�̰Z��u��qzܝy��l㭽f�g`Ɵ�I�9n���*)~�u�c��q�sXB5b�|�5��y�h=n�	��Rq��B&����`a���^�7)���� E��&���9a��|A�5��]XD�q��\ϖ�h���:�e�@��Z�N'?��4��`:ivqh���s��<,���KqC��Q2�S�K��pԄ�.�z�\�P5i ��z�G���$P�����y��^��_��,L*l�k��cX��o�N|�_��3��Fs�N��4�B��u!\e�������E�x�*noi���R�藰8i�E9 ���׮��1K�6I�֎�Z�0{����.-b���g�~�q�$�����!�����(�K_Ǩ��	�]�*7� �K!b�6A�$�e�[���)|H����+6�K�̈���!i�#��N1Q���$pS�T�Y2mI���k-��Ѭ��tW`y�ݵV<���x�kњw�@�iD�x�/	�f@�]�qi�Wtp<C�-��F�Z�$F._0qݘ��?�(��ƃ��aӣs�)�!z�DP�*�w_�w+�sڏ%g��7�	��B�:�������	���('qn7��i�^\�}��r�`7g�z�X�����k?������[�i�z�l��6�m��6�*����EPl	NW�#�s%�ELr-��Cy|z<�'g,��c������ih�/��I4��R��{�)I����m-Sm�Ӱl�U^���v����5�J��u:�B�_ߒ�릋�����bq΅�-�u��G:�dѾpz�QsGkc o��wD����I���1��j�����-��uf��n˘���*���P�_�w涛}2��IфI�N�.�'���{���#��N�?V(|���l&TU�����Q���]vң���E��س0�v1�x0M��2VHNB �i/�u�!B~JPN�.\y1SZf��
4rm72����5j]m��_���C80��_2��:�U:�Z�7����r(�h��3e��P�d��q�2SRX�S,�8�j�i8��P"<�	zzI��2:���t��֧N4��{��{TS���!�D��V�i.��DL�)���*�iV���E��џ�r��z�`�W�����Q׎�c��8`(r �~WP"(s�I��	�L�B���r��j�вg���9
�9 q��Ϸ�a����k��O���ʒ�:�������*�4�<'�^������Ҷ��ӭ�D���4�������zӫ(LNC�HƢ�ޓ?�60-q�nhZU��}ViH-@�}�K����A�kb`4�f�	w�q=\6S��4bB�-5��O[���y FZh�\K���������R�Q��������e�h������ڑ��)k
�ږx`1س�M��s�����u���嫏14���5M��>��;��35G�i=&�r5|��cƐ�i7��ű��� оS&���\�;h�0+		���/��c>�(�:ʹ�J�-�>K߫Θ ���ķ�C4��L�Ym� S��\$-�Z�8ُCU-�-JU1a�x	+�/=�t�#[>hiUU�4��-�-���Wɋ,��OD��M���^]���|;���n8�Q�!�=,��G� -���K��͸�E����!���P��(ob�����fI�ֱ�C��@bjt�5�ŭ�[oܝ"e�D�9�O'gRa~��ݹԑ[qo�>�nP/���U�vr��+ũ+~�z�F	�>�������cE�]CM�}0�ML�*�?�x
��c3p��Qo�P�N�V 2A$`�B��?t+�\7=��)��0��D��|�Pnk�����������Bȯk{�rG�%U/^�o[:<�Q>'�u���_9s�QX�ڵ�k�X�a
"��#�#}4�{.�ư(ƠfLFS%p�p���[�� iFZs�iocל����@���/��NV}��R�;�#�̈V�K�}�	�h����'Cn�B��v;�KIo�̌hϝ �@K������ <M�e_w!���o�|��.��o�Ds�t�(K� ��+.���Ԋ�O4&�3ء[�?�1��)r٦��?�a�R�myz���_-���DY~�
Qۅ%>�E]�$j5��+,�.
Xplp�1���OqJ3��[f[B��c%?-m���˻5��������]B�������Fn��q1A�� �=M�C\7�R�W�uj�g�w�f� w۪�0"HmX���P�ץ���$����q�~i2���8O�utB��d����k�n�%)��h/��ˑe`日����h�ɖ
C�)������.�f�Dy�ld���ڂ�0�B`���L��n�^�r�0)��,���#���K�+n����f��W�Od��"��[� ���Y|��^n)g�=���?�s�@zl�S�z�2:�Vm't�jN5S}�X*��.j��%�����v-{���n��tCH�V�)�W(�biߜ�h�7 ����	��d'���ޠ%�
���Cs��n�DJ���}���Q�&���
'�ވ��B�@<Q-���7��h�x�tN�6��,j�B�ȗc����R����FR�f`������Vuq�S:�x�*�&�9�v��t/UXOA
W��,$E�׻�m����[0G�۞�����n3Ss��b+�*�a�Qv�5��z�ay��!�Zd�E�W�ʇ���[�3,���o���l�m
9�=5����9*�,�@�̆Ţҏ�8]7�h�	$N�܇!e�Ĳ���=��C)���I��Y<���E3�����,Ĺ�T�1L������������j�����11��� �aZ����s#�s7�x5�@��g�'J����u�y.�0��"����tUʀ[IC����y-�'������IJݺ���4O+���j^�p���־���-��o�\<����dc*!%���"p)�ndW�p4]o��f:\�[r��,�ϱ9�����|>��z�G��T�޲��b��s`F%�H���"z滅JZU1�6S�%j5r^X�X^���D�վ`A@(���#X�����B�����BNF�n���5P����W�v�:�B��AQ�M���S�8�/�,�ș.Q���\�8�(�>+���ߦ���� �M���+�?D��bS�E|w������0�_2�lȒ���.$�Zn���_����`�o�3r�ξ���X|�	ja<�zg��ɠIH�ߞ�,�Ȩ#�K�%���Q˞��1�݇
qPt���$�j��&D���o�	����B�ӮH$HLǞ�%@�H0��H���)K�'%O-�N��������]��k^��DK�9��YȽ�0���+�b'x�/�H5�z��}1�$�(����|C4h��:a%~�fb����jt�e�gR�d�*�B�k�Ա����2ģZ� �w�ھ�.Ә�磁f����|�I�).�1q��6�'��t����5���'䦉��?�o�o&�3��9-�d<��Y �FF���8!��!���Iu���"�h��5 s�����oG#?����"�:��{D	ɀ!zԆ(Z��?�@T2��%䲜GbWH~���w�_�[(��o�آD�Cő
����Dy�g�	۳���h�l��b�Uj�{�Ss.�Ħ�Չ��E�ƽCQ'�kL�3;�nHG�H#UA*<S��G�մ#P���N��O> C$x��/n�X���̕F?�?Sk��2�$�����{��Ǝ�Sm� [�,��_��$�5�-�&>�E\M��g�{����I����-�V��^-�>~f�b�<	fk�$�ݔ�Q��LQ����R�����D�Zh�+e�S�Z���yn_趋���]��E<�NV�8���'�$5�y]&:��֌׾ޑp�\q�啌����CpVU�E�0*[F�0������Y�'� O��R��¡Z�>fN5+1�!�H�!������d�����ʧ��ǔ�M����dH�7�VA�@�A���2�c�Kӝ�ȣ�����c�,�iݳ�C�:�h���U�ͻiA�z���/.����K�������e�ػ>-�S�x��o��w�艀	�����:o_?���5��r��"��GX!�̶�|w���@��7ɑ'�ԧ�+[����-}�S5
ֻ��æ(�
�hkVZ���(�/�)) �vj��(�j�k)/-U��cfg�碎���3�^2�k��0��S�p(���V�c���P�#�YS��ox��ů[to��-ި��ޢ����SK6=Ƭ�Ӫ~�y�es�U��ڏ��c�3�%7"ؚ��K�W�����K��o�XF�'�v�'�LG:��1�Tת5�{�2H�@	�
6����a�� �T)r��ל�u�<Om��@��"����SnlUb��{��f����,!�rC��E�Ş�COZ���Ymt���)�[��훗u���$`��]�������������7�->�ӹ^fh���J����0��mg�}Z��lAP?��E��:%¤Q�J�7��ۜȊ^^���� �>�i-��2�әfX`������y�.s �sh��% ��v�r�CҪ��j^��P��������қ��`e�ŕ?�����jv���/�N����r
��T&�Z�M[ۋ�[��k�4F�ۢ��k�÷��v�U��jO��o��m��Px��1��ۥ!n�X�� .��.��̩ݚ�̄Q.߈a2q'!7��-?C�\U�]�.��!��r��<���!`o�Q�=J�2� B�{�R�(F�WdO-�#SX+��Ȕ��vy�P	�|#�U*	��*�Xw*�dc�#��ֱ�G�G�������C<���c���0��7��q�B
�>U	;I�I���݋�L�gM[��`}��8��J|�*�)h:r9���AΏ=�_��Z��-��V�`��g�gk����8n�J
����O.�(�+�/��Н��#@��4�wE��6�����A��W�����J����3T9����1��=��D�i5ְ�r�g=�p�����[O�ֺ�S㈠��rʲ�f�&��\� �e�n��F���&~��_; @�ceӵb�J��酑��7 ���v�������9��E��"���"N�qņ�c#K$���1��]Lͭ��'znphS]��N���0��5��qr���ϓ=+H����h[��ًC��6�O�o�{�KL6W|��0pe$�FR�O=�O��2�Ӧ��z�h÷��a�_&���ws�}���?�I�b��k�+��h�k_;��|l��;Ys��C�����{zM�&��3稫q2�3T��6J��Wл�Q.���Mi��	�J��;ԷrX��Q�]-�Z�Qk2��:�t,�O0܀p���������ǂ�K�g�l���?�I��_�D�r���l_c� ~v��H���[(�gqf��h���v4#�D�b�y��ΰ8���W��T6� ��OI�G$�d����K�KO�#(U�	��>���&���*�I�I\� !��J�e�t�����QSq<���^�SR�n��y.	�km� ��2����H�NbW��3�F4�=fr�{��,�o�O������<�w� �w2�+�zy���ڹ�@TJ�Q�/�K+Up��/
A�+'��8��$�0;),P���e��������B��Z[��F�e�`v�I��\\�:��t����փ��G����񼘧�8�c�&�unP�f#H���Φ4��$���K��ݍ]���-��3��@��B9o��־#��H���hOtz��f��Z�aI�_�v���;��e�+��4��PDr2��Zy�9��&r��cm$�H���)�}��"�F���C��n����w�n�֩P���1�c����C�G����ᆛ�/�R�P۴�p�(��<.���۞��1�^�V�<�p�v��7��Ͽ��ʄ�M��	A��g�M���J����,Y������j��!�|+@d9 �f�s��+!��m'Z<x^��9���'x`���$C������n�� hP�=}�sN@��koJO$��L�p��RKԣ/K�ey6�����I�H�����c9܅����`�o���hIvt\�{mo�$EL���2MC��s�C�W�?�;U�y{}�R�k�,[7�s5F�Vh��\tW{�H �~/7�Lj��vxC���5\�:�}�TΕ��[D�Hs�6�?�K�C�[��z��Ӷ^&S��� �p{��,(ZB�!��)���"�u��r"���Ab1t�J%U �Dq�����[�ΏT4g�0��d<Q�!�}�V���t��ʀbUjY2؞��5��ͯ�D��E���Q���sųVp�$z1�<j���O�R� �ӅJC=k�םtL�֒���?F0�K��wR�%���7"g�Ⱥ �ú�H���>��'f����:��2��?U:d��]i=���8W�kf�ɈM��$>�]��t���}���;�zc�Bd'~Y�R�b��o~�:0�%fx���44�XhFl�o� 3H/�����g�*H�E
jI+{�@	��W�	v7(>�[��`SF𝥣2�A �Uq�TC,ߤ��"L��U>���٤�V��+P���8v7�n���eWx
�DSux�QYm�rk팔u��d���y�o�m̤�	^oV��0��#h~Lm�l�<�{
�k7l5{;	w�%�����||U9>����7��O&u�zY��~��7ȧE��W�A��G̫H��s&��[tH�����
���g��$����<�g��z(�T����O16�I�qy��U�r���j1�Xn`/E�V�8��~=[�=$��-��:QKY"����
�M�r.����w�^���|2���y�}�G�-����ֻs$b5'��36K��yw�������p��"է̀-�<9�w�ogj��|�#v@�������ҧ�[L��"'���JS�qa8�ku���k��n�>�4��VU!��u����-	"$�&�ފ��cQ,؝���*�D�I�d�O��%�#�[f�x��㠯~�)t��bjO_�1_�3A )K��l�۶hn&E��%��������k����W�>k[�Vg9�>q/�ADzw�%+䜮É7�jv5�͇Bv2���PA�sM[��U��R���f*I���Ϸ�05#�~�Ne!_&�FT���x
:)���>��0y�@��PK������I�d ԳO��G��u�f�g�a�u�� '`��O�t�En=8w�U�F���)�x�
	�\��Ψ�,��F�6@�t���ݍ�]�D�\��*��9��u��� Uo�cR҉r��=�:иcˡE���t�>�;�-�A|u�����<��t����N�Vۼ�E�:iY�*���%�p��A^ӿf�Sq�D��<+��%`.�ہc�<���/}W���p�<m-�gcn��p��3�>���5߀z�u!�~�.��T�8�[gV,#z�q�����r��r�1uyoTuP��:��锧�J�o��Q�q�>��Pឦ�LtE>q����J�����'�5+�#��	�th	q� �Kb�ņ2;�&����yz*�f��7rF��tE!�?�N����+������0�����R�T���X(H�4�3TПB8����*l��������$|�h�(�\d����yx���;��/�;����ˏ4V�=�}�8��0ZX;�N�vW��.-顠�����0oC���+��	艔ݬ�� ��Q2� -[��G�OOПE�0�c_nD��b��al���e�s�L��¹i��XnH�O�
}�U ��ל�"L<c�����*�{Q���=��m�]Q	�R�.���D�#4p�W�ѬB�4�O4��S8:1�T?�he�Y�"�����@f�+SB
���ü�#�����'���y���0O$n�D]k
�H������Pp��!iN��]����fH�As��{�)J��Po��jdNֳI-�tM�]y�ע�;�&��ũ�<����c�5gi��G(�=�����~�k�O"��$}����H-��`�7s�ޫ�Cmpx%��9˫�&�������c;�(/�گ��O��:��L���94�0�Bl+���. ���WŪ�?�[��8���na0÷T��֭j*�5FV34�O�v����^@���N�a��Ӯ����w��5��Z�㜮��ms�c����$F���5�5u��Ľ���L-2��~;��TXB�H{�����S�� ~"q� ��3K��V(ȣ�:ĺ�pb��[�O������u�:l�-�:�k_���B��{�3C%����	���@C,]G<�]���꒶����:ty�Oم%Ӑ�Z�%�D
Zi��No���8���<�/ZDX�U'y��Y����--L�W��[��%ؗ��(6*��+A�4�H���2w��-��O�g�!�3<}܌��&�T4؅5޸G?W��ǈ�_��I����]�@9��*LC�