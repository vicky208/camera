��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G�2��0m[E*
�*p%~�S;k����7��&@���c�q+#�$�[$���gE�:7��P7��X�3�~rq���JY�#�7�m���,\�|@�\'�����P���a���U���x�"�}�{���F�J��	��!m+�F.�2U�/7�v^b�jI@�80������u^�}a�ǿ)�D�@�[�����J���%����v�Z��'�ļW�mr�
)޵2.���9'�FQ��ҋ�H%+E5f�9�F�(��C�Z���}�]�>�I����Aѵ!/Dm]wڵS�C���8o��)��M�Gi0���y����o��]���f����h��Z�~}���{��|'a�	/54`}o�D�$��;#�ӄ�E�9���Ft�4�"쒋����
#���{���8�������|�}$MZ�.��� �R����=���3���������w�_]zm���h�K����ig�������#"��k��X�����e�z��d���c�����"9k�"��E��>�^F�d����]ac^��I�K�=��B	W���<���{���)o��d��DI|������10���b�W��Ȝ�tF;9Ϟ3�.V`?�e�0 6I����l^m5{{��׌z��|�=�66����r�
6J��uB��8�+���h���V�/� =��$�����eu�Jl��\,g�a݋9�Y�)+��\̤�e�?���w/6[.��[]Hll��'J^��s��V�uc��;d _Ch� �7��6�Cs!S���Å5F�6I��K�]J-�0�|��E�g��8��7i V�A,�/�z�=7��@�f��4����Y�J���Ù�W]Rw�E[wT��`I^��zV��gߎ�ϱA t�Gq�˕.�8`�9�Kt�Ė�߭�Wp��n� 	�U������c ��-gyҴomD��8/�W�H�آ�[����\�%9��C0��:��е��
��jX�J_
�k���!��]Ї����#l�}$����
�eh�Әo5��43���Fh����<���T
P7�ÚvLT��8�N��>���ؽ�]��.���hb���╁�7آ*��̨��j`Q�P�5+�%Z�2��)M���Ȟ���@J�M���Xl�e��[��wß����3y� ��cL�R����h�d�!`�;�S|���(L��\��I\D7~$ :�P�4�*�4ij�V�@;��
Ô�u��'��U�������,x/~��!�V����AA§����R�i@��H�:�޻+��h�D��-s����e~(��}=� ��#��$��
��2�M��%$2=��k*IU�s{I?�����9�s~kqj8�fMƃ��V΅�a�y�͵�j!Y�l�qJ$�b$p���׿�)��.e�n7i8� N�%!�en2����*��>�AJ�%��>���nź�0C(��4P5@p6 n m<:˚��+���&Y%vM�b���z��W��NĭX���< ޴w>+��kF�� ��&ߧD���J���)y#���!'�=q��}A{�~B�?c�e|�)�j~��o'��j�oOAhW)"[c�m���9=~ ؤ���-�k��<3}9 �4RZx���,1s�Œ�WO�z�	Iƍ���[r�5H`��
��/j6C�9zK�ݗ����O3�&V���f����ñZ]xA�����j�>�u'�D��U��*WϪL���1�Ӿ1%�"pv���tJ%�� ����F+�0�|�����d��O����?��Kn�"4�1��wOGa����Nm��@ᾑ�Px�3��2�O7�!'s���Gnv~�� ü�8R���O����T�џ܃	��R�ʭ��"�d��VOt�"=^�E"��Տ�T���<�,$���g��>ɲ&��pϳ�N[{G�����w}զN�w"$pk5�PA�[e��?��i���@CQl�A%���-gl�<7/���Tg{\=��]��Jɠ�	�O��M�(��O	�Q
z>U��f�tH��m�'>��@>�R�Mn�E��(R�/��Ԍb���7o���Y�,T_��P޼mM�{RK�:/�kC��V'&���U(�I&m{�k9�ɚg�<�yAI(VD�	�h���\;�b�z0���-a��Iq&�C,�sU��F�E�QS���u�s����yT��YA_�4!�L�&v�GK,��D�`��	-s�\�Y�_kT�
�i��s��Y�V�sS��n18��p�>U�J5z��R���=k�� �_��A l-on�1򼇻�M+������_�p�L�!�\%$����NvP��6�R��/ ��T-2�~�d1�/?�$j��=u��(�����F8W�Sz��L꾍��x�1�Գc��+����W����'0	��e�vO|s��4��k�.'&���F��_f;[�S�P�p�c�Ş1�U��l���'k*U���]�b?N��Ӿ5�d���6��g�~��f��*���KH�2��$����Uv)y�i��ּ+9Y'���z�@^�j���J�p�P7��!�{uL`�5���  ��g�1b�ea^�`��(��*�T����P��֥Ȇ�Oq�#�m��.�Ct��?�O ���e�1�{C|$M���r3f���T	�]�k
&O�RlW�����e�􊕝>�'�ٳ(��6MD�3?Uk�Ղ�����(~ҙ��& x�c�n�p4�+U��;4 5����V�;:3k�Ƨ��-n�%w�g��	���;Y�ٌ���qX#�GQI�nŁ��z��o���P�vB#ȃ!ڸ*
����m~Tc� O�ۧ72c�?[��<9j�d�����.�b�q�O�ᬞzo��s�#
*����;��٠%�6�Z���|0a��l���u1ǳ@���n/�q��Z�{"B��Y�'��;��-V�$H��ő��������uO�%|�"�֔>4�]�Fa��hx� ������:[Wʬր�!�:���^��Μ�����Kuo��oԝ[�:�A>
M[�̵��\�4)rl����m�B�2��wß�������P�HY�U���a"�M�	x�g�2EBR7��"��bh�V��I�Zof'M�ȧo`b<��M'��z^Mt��c�<4��?	�*'1�/ 
,w�9�.-S
�M
��x���ۍѨ��c)��eg�����<�~IC�W�U�:����UH,��7�K���n�[��Yp`16x�n氝��]��>�غ��?��@/MIn���%��ޫ�jq���&x'�����Dm:�-AXd �ʝ(	�h�QZ$C/'#_�kR�Ʒ�s�5���e�6\C٩�����>}~��,~=He��L�dNC3�'������ ��ɱ�4|��v�7d9��	�[t]v��:����'���lY2ا�_ͭ�b���*��.Օz� ZB�s?1s�PL*���1('�p ���v���9Ƙ��܋~Y)�#ƃ�Gil������k"��2}����!���5�}�)�ŚG#����_�)$��=��q��n�g;$MO��nh\��7�a��{���j2��VzM1b�c�dӝ�\�{�.����8V�J~rH�t3}Γ�cp�.��B��,��,����-i�[��g�=:���������JH�)��˜X����"�*e��f�LՅR���ƨ����cFt<!�=����TĎM���tfk.�ix �'龂�1ngo`�N�}�0����6~V��wUY��z�`Ā�"���R�0B#O�#G­���1�%�l�8�Q4x\h�l<�ժN�<MM�5-�'�w�O9N��y:'�1��ER�Z�ۋ^������)�	���O ������$vo��1:wbԩ�!D����/���ɤnց�E�����W�;��}&�I�_-��C�ņ�fG�>>�C`RZ��Z0�ߣX4��6���J���6:��mH���j������'�����sa׋O�t����W��s��.n�3D0V�Y'���1�o7Xj�~�N�5��f�Sv��g���������DIF�7��6��~�1j�P�=�࢒4��_�������'��$�<&�O�yl(G'K�4�*5����ُ�8HP�4��� �=}�&mn��0_�Q.B��6�_X.�K=p�6��ܬ7�[�w`K}�[�2U������,.ro�
4��,��i�>����������-�[t����p�F��|��`��A��*\��#d��mB7���C�)�94����J�yh\�>b� ��K7/�E�}��łNz~�aHƘq�yW,o��_��x�1�`MR�9sIBv¤~���jI��9q���18�o$�ꭇ:�x�Z6�H����H���q���ߺdx�p�I�K)� ��|�y�/es��?Ϭ�d���5C��m�ϡv�$CIۍ���E�c��J�{AD	?�1!u�t~8��)P���#��ӥ;���q"�9��M?�V�n)��x�l�Z���73��RЂ\�x j^�^?"���i1�!����<	T�ùMf"��]g�:�rG�xǒӵ7�����ԟXQN��u`Z���NEJ�S�=GCk�^�����W�t#�pwQ���̣�F�]�pl�bxք�w	m�=~�̖�ͺ���.;`i&\ żOd��ū ��TU�M������Z��u`�g�(˥$��L#Ev;k�;����o� V��rۍ=j];����3Xz�������*����~�$�<,�1�y�몏��K,�ӏ�&��c�g#^	�%^�� �Z��φf*�[qy���z'�kV��(�|n٩�VOϿee^����5%�VP ��	���<�_����6�ɶ0��E���5��TI��'�:un4��Mv+� ���������,��
� /#�+�pr�.�x�Ҡ�vX�ߊ��^�Iu�N	=���X����ҎB&m����<8���7�Ɛ� ����F�)�v��=%R�;x�HH����Ŷ�E�ͪ-῞e�νA~a[ч����L��ݱz�I��:+��8��%�(������0!�J���E/�Y�J�݀����$��W��j�a9i��n�N���u��ӈ���������J'��^�@ș��=�I��DXQ;�g��zQx�#�$��{���ODne�5��ڴĶ=�1U8�5ٲ&Q�>��x����P"V8DAf<=�G������5z*��R�����6��[י���^}���5�eo�=,wk�z��'�3W���'f����)���C�S˫t-a�SA�_�W�i}�t�{��oW�Z����"dZnM����w��n��.\�5<5O`EX��6�r>w�UXB\#]�ad9����'4d���q��쑼$������Ȱ���Dg+��2N�zI��yʐ�ͦ��&O�9˶|�d�y.�+qBdayMi�*����8����'{M�>4�x�g=	,yK,f�pU|����x~�o��gW��ZK2���]F���t�{�(N
v�ʻ��&������6i$X�"�H�vlw��S4n�T�gY��4�i�	ʍ���P��X�����B���p� ��[�U�H���~0����\��U����
��OeK�Rj&��oJj�v��{^������Ey���c�	P��)���\|x<�rS�|�U�7R��Go<$�u�M�O��q�)���@�pz6/[��wRB=H3��~Ћᚐ}���^�u��7�=��i�Q6Q:w�s��	��������Q�3��7S!K��R@X^��VʧO_���V
�w�d��5v�qʫ�����q%OM<:y"*\���1ߌ�b��{����0֯;�l�"4�ON��9��	b ;���Kl�ƃvd�>����Y����� pQ!qz-ˉ�U{���@��<��ϫ�����4)Ưɝ9O��p8'|8X���0�&+W&-n���}DMz̵Y3�E�?E��4�N�'v��a.���흚ݿ)H��b�߰�<��<)�����M�����t�0��r��o��(��>-�T��<�ѯ
Gŝ��O�iz(Mϥ��C�������J��+D�M<	.ИQD���!�
�؄)�xaX��bW��\~PXP�榣\�3�>���o�u]���97A'�}e�������3�s�%�}�S*io�)��Zƃ�<���8���n8C����EM��w��j����T��#����Z.Y�5�>���������9�H�X���@��x1i�7ݛ9�L����� Il���QǓ�{�E��0P��]NJ�G�H?gJ߱�?A�Zb��6"A뚠�e5�(�m9�×"���/��� �ވ�� X�uQ�`
�W�9�w�	�
�y`7�����pW	�o�A$�m{�گF�ޥ׌���zY���/�{4䘃ᚶ��_�+�?������p�Er��Š��P:7�n����>�!a�4�Ș9H��Q ��Z�F$�=O���<U�8����<4�����)i�%��tj�V"y\��gyW�j�S
���D��f��[����%�㒧7+|���� {��֏��HP�Ѽһ�S���T��T�61�(Z�t�7��~p���X�]M��S��s~��Z<3��3���A#�8�N]�����A9l�w\���*I���ʆ��������hд�������U"-��r�D>���^>��>B?�d��\Pˢ_Sj�J�Q�{hֶ��x ��T=
?_X�!�N�+ ��N��/��R�8t�7�J�A@SQ��2@�px��ʃ!3��S�Ң���z�z������<���n+�T2׌��;�Y���l��Hov��Pw�Pt)�xj�� �m�RA͎: p|	i�i[�5*�"�8Q�΢E�t�s�t��<���̤���EYr��U���_v��0������m},3�f�us�O�Uw8�k��*�1�;,Q�0�XF����0sqB?'cS5�hz��_��s��5��l�'bdVsZ;$8B�>Q�F���d7�d�e�.:LO�]K�o����@�>uGr �p�[�a?����7r\]#��Ͳ�n�U�����>B�sVڎ�G�C֎M'(`��	Bz�|	�����̠�V�l�z!�%�U?���&Q��1�;"b��O�t����I�	��OtPSm5͓�2����p?����(Xc�J���(����ch���u����E���p�έ[~����4n��}��aw�0e�:�������.�r�y�f��w+��QA���oF[O:�ͮ�Bej@,Ǡ���4�xp� �8��}��.� �,�	�C W�ϗ� ��XL%F�Y_t͎���G�R���C��k��prx�
?��9)8�8!�*�(%A�}ڗ�1�F2�� oQǚi��!�%�2�Ág ��#��E݊#65Zս�����t���c+˳�SU�A�QW����t\�	gH2P�r�2�ByWî���:���l#��&�h:����C����*a2�}%��.���ו|��/g%K��I��;�9�h)����jV��Kzuq-2�G�/�k�����QmI����qs��|�dCʫި$�[ǐ�\$��1���fc���\Cz�H%a7�?G�@��_.(�J��[�!�ʹ��v�YT�� �����䕒�0���j�$�N}��;�1�4�WO@6)��x�Ц/�h�2�;Y�8c�5����aR�/����6C��-��#/'��?tL���ƾ:��lQBi�ح���dGxm�Jܽef���j�������P�� v]�Uu��\A�!�=󷼅�����2��b�	�A���r�A��]	)n3%��H���\�s<�"��n��!*l4$ꚞcJ&���L����u�����"b���R����>�i�H�gQ�t�VM5�vE�<$_W}���"�.���5�f2��}3��r���)�촨E?�b��K���S���.�[	��ԇ�����F)W�Q�_����4���3�����b[����r�m�@o�d�)�t��ߟ���&I:��l��6J�SAM}��UVT~�Q� �ř)p	���Ơ�߻
��@G*-�,T��ς���g��G�)��ک6=ӕ�|�����B2�Z���{w�Q�� �*V�����2��8z��#�azT`fp�7�|���X��<�j���V/�
0!(�K����9�k8��ܹai�w�ez% ���z������B�63aAD�S�,hJG�1�@�űl��>Pa����"\ǽ����(n��4ޏ@��~8�N�-
�<Í��y/R���7.�&�=�����I͛���-� ��T���*�"����+�#�>�Nw���%½T"�e�R�k]ڳ��4���T��I
]%D��8t��)/C3g�����Y�\�;|)�R���q��@�NO��+(���tc��wa{�,��$J͗:̟��?.+�E�1ɼ�E����v��C�ED�}�֮g�K��cx	4ױܢ�p�0{ɶ����,a��������&���M�Q�������S4�ɇ�����]{���� y�k��J�W� 4B��)��?��� �8�������'��!�!�Z�Y�n�&'�){�/ �f�f���K�7��W�/�8�%Ӛ��p����GWw_��?'�@��s(�!Bb���>DF�c�mO#���O��c��H���%����L�j~�X��U#��7�R�����D=8���Z���^����N�#��ɽ�9����px�p }R��s���4��C0n����>K8�#��~7
���=],��#�9Y�{�1����@KMmJkG��we�p`��������|y���}ǖ���6����6e�H�ٟ́$���ܿ��-8\h��x�h�����\����	���_�ayB�A����Y����= Qxm&_��	g�BKMXrVHq����&��T"G���e{q��.#֏�R�����kȶ�<�����b=�}H�S�*���B��}��I��͋�	!�]��y|��aY�5㵮#o�_'��3�%ro�Q�V��U� 4q�Sz����q�k��)5�	8=p��ʑ��[zH_
uE=�}�*�M�SU�A�޺��_�m�HM���ţN����-
I���7��yj�_��k�l/�iM�)���t9p�T��a��4Ϻ�0;dH{�:ڃ2�5:3Ta@�hH��0���>��]���z$\�Wƹ��햗�����N7Ir��ݸ�w=�:�F�����K���!3�	V��҇���M��C���s��V��{����<K��=4 g���7�Pco�ͯ�L����q;�>�� ����i���t�Z�c�����`�������d��N�^g�x��pk����G���x�8'���ҴU��L~x��ރ���U��~⽋���;�z�$�>2�R�*�����DWwST!�0E��Na�,�D����6����\���X�]7����3W���c�&�!{pj�N+,b|��-l�l��{�#ә8\��,}t��=��"~�r���j�/��s������22M#��Xڹ6�����<�Z7���:�d*��+���G��\�1z�e%��K!���{|b��8��+ �A�]�&�F�,���*�.l�LO1�V	З��kv��(J�����: fr)OƜNYK����aX��ݳ���5a}-�P��g>���@`�MR]��V�����f�N��"q�H����pU	h]����l�g?pZRk����%,�yޥ��ڍ�/#��e2:_��#'�i��v�p�:&L�\�Z1]� ������RL��q���E����TG/G��G� n�kgxn���\��S�+����������)ϬN�cUg�6��2ղť�1̤Ф�H^�C �Y ׁ�JI	~ч�Wdqa�R'��������A܅M�+M-�/B�K+�އ�QJ�Hns��y�:L����BXA����\�v�wQ%�}�;T����,N���4t?�)�J�[%Wo@2/��>σ��f�q�{�{&G+�@�SY'W��VA�v�S�B��t�0���#��b�Cq��јl t�\Mpn*R�����W^"�a=?ms�GmP�~NH�J���8k�	QP�F�*���u� �3�j@����/����j����4C��h�A�	�w	h]z�CJ���2tnQ�߯Uc��(ŷ��)�a:a����w+[�$��r�TM��,��u�����+�������R+W$1��%&�D���kp���p��4ߦ�V�"9a���7���se��D�S�!����d),�7�¯�d�1&-[
.��S6Ax���+�@�ɭ䤉��Ձ5���K� ���Ɏ�#'&��$xx��5�fik[�	��H�!y_����Ⓚ'����2젠w~{^���9��ȫ����v�3M��uo�	��R��	�Z�>e[w�[����F3�,7�����Q �X���.�4v��v�2��ޱ�>�T�����|��k�r�to3�b=,)׸����ǖ�7�au���1�駮%p�ګ��PC��
�: ���='Hc�Uj$2����P�s�zGR�����S���%�0�p���+[P�l'��16㻒�H80f��ϽWaKNx���� ������A8re�2���c�i�����l�a:;�5�Xb_VFK`�jլ�Y���gG��PE�sԣxu�^����B�?G.��lG+�R�_�6���P�s�:q�A+N5��x�±�/����c������gv`�r���I4���xޥ>1�j�I"��m\y��u(f6F�ӵ�5�1T����PA���^�oF��YC�%�����Ɏ����k8������µ��⫸��q�:.��8�~�O܉n�E��'��`@;�M|�$d=GrV����%Cxx�'��X{K���R�i:�ƀ<�ݦqK�D�.���PYb;b1K�I��!DN؏��֒3"GnR�<`+éy*��߆��3hO[����|P����д�w���S[��p�E=LR��M��+N-���_BL�ʺ��k/�Ml���i�4�M�p���HO-q��j�P3�V�%ke�>,`�'{��2diD����#f��t�E��h��1;.��>C��냋O�#9���hQ9$ޟ���vJGE�+�C~5,�
U/�gl��}��)����F�@�t�'�a�1�^�1nKX����rV��?���@% @Lv2P��Ƕh�v��+��	G �5(&w�ؙ��`�2Y�G�=D`�8HƉ����T9�0)݋	����jD����3"eTv�H/!?��O��3)�r�I���۸��<�_����P>:f�$�EA#t4刬���	������阭�m}�M�0
>�������E_��X@<������~Kq������c:`	
�Nax6��ȁ)�V'��4��cL��Ǩ�]��oI�����!�{.Hi��5�\��)��d�Iv�("+�Y�T˲��P�Q��=�)W��#O����@��5��!�S����f�ޑF};�k��8Wy�dX�'��gV�4�x�����	o���3da���l����f��������=�#J�.b*���K<鱙D!$ 1��9�����o��%J����HNu�/eQ�2��k��{7odgL�č���rE>��I�Z��g�����)���Ɏ׵4G���g�=�jЀJ������R�m�k_����[i��n�F��н�2���*ugϚ���\*XRM����GM�G9��C�cFg���V�Ds� �	���P��ʤ	OA��4��|OD��}��'5��#V"K M�;��(ΗA�+�p��Z��l��4���s� 'U���zr�rR����e+�A��C'��X��xt���&�b!$�6�|dm-O%	C��x�Ѧ'P���7��rN��|��v�x*�x�]�U���{jKM��;JH����C����%�G�E�� n!Z��4Q�&�:Ji�� �e��εX����D�o�b�}F��K4wޟ�:7y�V��uIvJ�l�27�MN�QM� ��@V��`��1�>��{��f�s�S�BR%��	N6���ʄbU���ӝ �����{|�% ѫ�[�.��5V��v@�|����U�b!%�Dl���L��	��@�w��۳�L1{��P)�(�ۑǛ�}�VWR"e-M��_q*p�3G�:�t���j4�����~O�|�%��K5��w=�Сi~z�^�`��ۃ�Z}�롞9��T�n�X�I���R�O��p�^�QT��O�����o[����-�,��w��H@�>�T�NU͒��o�>��
��@�A��T�,�w+�.�k��-6���&P�?c�q�9l?1���Z�>D�C��o�z�3����W=�?�&��g�O+\��B�|�f�
QÚ�F�pi���(JFpϙE�D�+�Z̽"��s=���������`��d��z�C~�.`&�G+���q4C��$a�-%�~��ck�Y�(��)E�|}�..Eȉ��a\�����k�����f�j�,�X:�י����p:��7�����/��dvar�"�D���`>�X��;�L�t8ЛC/W�$�:�~\�J�7D�� ��)|7�_���]�z�_�7F��F��fh��VƖа��Wg�-�uE=Gǝ�c��X��S��;ùU=3.����~:si�:�g-0�JnK�◩ e5$g�.�ȿ�N�E��|:\�-��Ƿ��ba�Lp���f�X[-�Y���k�w`�^�y�E�I�.@����{���u�Ʒ5��"MiE�]׼z�[��KM����o�8ti��xV���QQ�X���ݍG����;׮���*�rB�k����{*�6CK�u�c!^�����S7�*p 5.c���ݰ]�`8��#�9:��CD�
{=�1���+��d�	t���G5<�+G����� @�qo���;����T �p�1����pv9��;rb�g�76����%�qS����N۾��G�;͡~B���{Y$!%�U�DB��RyB�Ⱥ��ۡ�p��"��\ė%��9�Mú��[��G��:)~Xj.顨�S�V���̝���|pI(����	Bp}�$�Q&2\]tc\�*�6��Azn?ՃC��C��w�\������o�^�e.�s}Lr1GQT���W	�LW��j�^��"�4���n��S���� ~����#��t�V�K��D����R案/��Jv��lwR����8����?@jq��S ����[*��[0�|�zxD�����m�Ԯs���*C4��F���f��O��w`r�O��� e�ј��
g��|�{�}���k��* �z�)]�Pn�X	F�λ���xJ��h�0#!(�:g��8��?�;y��r�g*3���}��aM����#W8`��6�6Q��>�(U�hח3�W�IH:yH�;�hڐ�*i����_ԣ���0�E��*�~���@�"%�o���k@	:��v�pi��5�� ��[05}ҞF�f�k�\P��Я1w{TX�]�Iq]x��O���:�fdm�Tܡ:��$�&�48^c	�|r�~uV��-��?�VG���=�`D@䁤�}��3�l�>ɘ[����7`L(����S���e���jc&b��g0�$���X���qk!N��uG���&�d~m�h�0��s��rv�f�������'�!�&(:����*��4+����=څT���0�O�ƾ&�yI��d�G��Vx�bX���t=�cO�g[�.�~���L�D&(�#�;�����|ط}_V0q`�k	&�:z͡=3z�%R���uO�f;���c冸[U���53����Ь��6kRЙ}��Km9@-�s��`X9�ɸγ�XFb�)�g���~�y��<Z=\��P���i� �#r���^j!T��"B|KPjy���Cq�[{*�X[��z]���R��a���'���F��w[]�"W���^�5U��_�_ Hl�b���z��C(n�@�@���	������z�6�Dz�����bP������5���4��d�lZ������n�t�U�@�>��A���P!;ȧh�C�IA��Ʒv�y'�~ߔQ;�2;:��ۮ7��z���ۚ�s�`�EC�H��V�s߽J�mw��%� ��Dx��NK ��s�~�dX��L�n2�S��7N��m��H���h�x|�g�f;B����܉BXP����{��n�-�5��h���T�SH2��.{#�Q��X��&��sr��M��n��I���^�d��KR��C8�bo��: v�_��i?�C}��b��3��T=.um�B�,�($"�2<��Fzl&0,�Ya��H�g���������g�?��o��<��z�L�!��3�C0����ZO>X�k���b5���ﻗ�8Y��[��7����N6����LA@��{t/[:����q�\�1[c�6�*���m�N�s��\V>Cml�+�3W�n�Q7�Kp�+�|4���.�6�?p�!�+�*<�0�F^�� 4(;K'�����e��X�ꨙ�Ji��-��)�,������PK�\+��h���P���)�ơ�!�Q7@F};�WmPf��ht��Bf$a�iE��?����^����;D|>���`�ⶤϸ�����Ge�@�c�d��B�B� ,����F�52��}�!��6��8%/��_���fp�ߪ�H���7���=��:ٍZ��r-X`R�<��³7n%!��n`1�a�ж��L�����OL@IU�����'T��m�t涧o�:��<�ٷ5_�ߐ'�|+��fA�z�	o-f��/���ի�.kI�$l�\�b\es�oI��;C$So��lhz|�
|�>j�/e�.�X��H�B��HG�-)�r�]4*X6��D.S!�`��߅]d�̈C���w�6����6A��_�i�}�����z�<�k"�H�5�8Z=���4 ���2yb�FA~��b�Ō����:K&�3~�S�Yd�`?�6h5Sx���1��1��"�����y-��n�'X<�8�O ����|J,u��nc#����gD���؁��mV"�A��bm��������A��~�|���ҏ%�S��6�s�a�O�IA[�sD.;Y��dys����Hٹ�u0��`b�AR o>����_��T�R�����
ހ4/�Vs�d4#;?9��_Xbf�s��2G5FH��'��F^�������p����C�T������~���\�B]xqt���C��-?@OD�[�dSa�P��c濳4��:�{�(�FA/s�`�����q)j8s�w�sg��"Hx.�ٻ>�B嬘5)�\XDn-u�`�I���dw�����Ce�zj��9�x�R�2��m�=���jh�[��{҅���,�D���!�g��!g�ڸ�"U�q2���D��� �Kw@�6,t@��J��(��u�9�3ZL� Y6��$��]g�9mAfz��	R��ɷ���>���ǎ�3,Ϸ�p0kx��P��AE\��l��_�r�H[R��N딶�^�����-��>���e�U�Li.��8�^��0�բ����G,�Þ���ܕ1���C (��YC�d.N<��<(&�G��	FG����
��)0�y�~�+ڷ�ɋU(+ˆ���$��,pe��uE�Es�z����Իdٮ�G�Gw�6x�ǭ�8}�|�lc�t���A��t��x�1iw��E6��狈o��ͱ�>�o*����);��fn�!�&	�E֞�~�ى�M�f�; ������g�k��o�Ԃѐ,~�W eA>����������0ɦ�@����O���=��ө	2cdmF�`��xPS�!T���c3.�/#Ya����Z���[���;�������d�Up�@4�w"��p"�#�䦙J1��t�K�Yr\�h)[������#qj"�w&ڞ^B�Ea���U�B�kԿ��@�����F�_!��9��u�_�iC���	 ���Y�T� �8��4l��v�]27k�S0���gar�Nѥ��y|��[��%`���=��i���7�8س��>���ly`6��{��b9�e�sE�v���fѱ)���n�Ft{���sY���wW #�)qũ�,'mc0�G�%q�RK�g����Ob����A�y�8~ɷ��c'8'���������~8{Zϛ ˌ<XN�Iy��$�?�����DC&u��پj�u��V�Od���fgkF�j�urR+d�DU%		Z�om��4�s���m����W���c�� L_�o��0�䶌ٕ���J[KTZ�����j�� �g�Dxef���\q�����O�|ߍ@S��a`���	�D�2D"��8��(�u���P$C�6Q	\�����'\f��
r�����N{?�����jE� /A�jf�m氖hc>��{�s�*��.K�Z,������T+��`�bߤ��r���}I�P���聳��cKd���]a��Xۚ.����C	U �����'O"�&�4�8���+�T8������Ts�1�$g���o\bci�0��eA�����@<�y�28�v�|Z�\�	�Slv���3���&�H���SB�)�9�K��2O��ʣ�{�{�$���	�T�ca}��T�ӎ�T-�q��^o�ԭ���P9���^��1��W��� �}���IY�*H.i_`�	�ʓ��.cL���N�V�G3���mӸ�$/;����r�cXw�=6��f~�X;>C*�.�?w��!������o����C{���@(z�C��3�G�H�@�t]+Ea3v��K
]O���$��d�h��?e�KV1�}�	���4��Z)#�@eюӇKo����P�����\�yιM8�R�������pB�z�;��	���YY�oD�o`:�j���f���$��z+V�P��aX#��L��}춮�w��+�4�,;1r���?�>���G܆�zQ�
�6y�=�z�]�Ѹ �]���d�Ǉ����,�\{��#f��[��>�Hv8tK���啵�4�5^\d+Y��/q��#dr��ۢ�>S�Ƒ(��q��E��h=�LwY����\-���b��?�v�ȍB�~�؇}C�L��>�;D`Euf�P����]�{�f�p6ϭR,��q�����NS���ś�ʒ�PA��H�j�L��}���H���3\a]v2HIh�=XU
W����w7�긒�L\��31;O���������w�A���+f��L�n��T��cv��=������<��ՠ�M.};죮;�:�5:�9�f�5�O<^�	tY;{��29ga��(m"�>po'�(�R�bΨmP6���*>�>m������,�]PE
KŘ㙡��G������^�0rN>���C`{XF$!2�p�7�E/�k�WX��[��nb�aK����-�� ��A}M�\)j�,��o��o��v*��^����V�^�s�Kԃ�R��ј�l@6�7���з^9҂Q����#�����1)R�֗�c�{�Bi�F��S9al����`r���8�2��A���"�b����$_���qS��`����e�G��u�?��Q)�+7�I?�ƈ��<�[c��j���z�K�a�ϋ|������Vw������½)�k���PUn1B�"��Yt^6~�k���ä^P(��c	P��0�%�B�l��uo�}O�l7|0K��z�|��H!��gߧ��A�	�	M0�����Gt�h�#o�칯�?�o���ҦsO�����R-���n,w-�"��@�4����Ab����!agZF	��]�~	��#�-МV� "�L��"��d����dI�#�%`GBf��x��I[� 0����嫡�}�L6��<���؁�#�9�:c�%�wy������	���k�3(N��6�h.��*�$	���*D��`�������I���Y�{w)�d�ѻ���`���ȘrJđ�;� <|�vNKI���lA��A��p���~�>��XO�t�U;mL�i�#r���o��H쐇L�� ��n�����Кa�:^^�N��A�R�_Cپ����|>�b��`��ۤ.�R� G������m��AM���Ћ
�	�&�;�H��U����E�X X6./�4Kq>��<�}4��o>�l)I�ʧ~��7��w�b��T�U�yj_��������+�e�\J���Ӎ��X޳�*n��˰�%�6f��p���-����o�tU�AP�R�u9�"�z{��1�h�Y�ԝ�g�D��/�c�p�*Lwj���a?V�x��xF�7Vh�H`��?w�c;��H����>�M���6VR���ov'La���ő0���i��;"����M���kZk��z�����;��h�9���Y���ˢE�#�\�V#t�u����[�E��A�ô"�~�Sө���yz� F8.���]4��HVP��9Cݳ��2K�}z���7pќ ��g]�c����b��46�ʁ���  б��LtY���OE��xJLM��`�q�RM��=��EM��z��е���ʚ�Ɲj��@[�H<��������zj�䡱���t�}3z#�cy[���_>�o��o��V1;ӉE������
�fm��.`�x/Q��$���=!o1�tFbs1n�Q璜��e��^&xj�:�p�QR?
t%+���!?K�_<��T�G�f�7�� }��B}�z�ط����A\��[��.�`���b���<g����M� �G7�2�N����=jOD���oE�������A.�����9����0Z�0.ձƷ�=�r߇g�y&�r��iWU��9��x`�Z�)e���~���"ݢE��`���H�+BꡰC���c�y�~�Y�%��r^'�/��~�����2�;���b�ծQ`�50��ݗ��&�]��0{.�j��1)fsNsbƄ�M�K��qb�Ж����wI�����0�,`;��Y*�֜ �����R�	���z*W �6��̓����j|�3o�حl���C��Rj�2�w]��Aot�+�ӓ��@،�z>)G��Y,��z�������� ��.Wxe��@��Cx	+�H�N�xɼ��LNr���$�P��eA�Қ5h��(����I�N�1���Z!'���>al�3G��� �SW��qg���G�6Xl�AX��;u�� C�ԋ�28v��ͭA�H�}À��[�o��R@��W��.�EW��l�Mڦ��ͦ�QA?G���|�[<��H]����"�z��Vh�����1^U@��G��-iAT��yjC��H��L>*�ġӶJ \�O��/Lfw�):yT�}���hn�]J<C�r"�lq�O�*wB
�)�iY��(�K`�[.����h�*�{�}��q��Œ����������]p��wű�`��1��I�w�u/]Tl �zy����c4C�fr�ܧ���G<�*o�����������~�`ٻ�^�ݰXל�u� }���(�˝$��4ɸ��_�m�D1�*}�{�ښ����}9Ϊ�����R/�ai=!���-�#[�C�@+��n�´���i���f��^�=f�gt�oΝ+�f�(/DiF�ň�1�Ф���d|�M]9,3:���(����V+a��ߕW-by�B����H	�6="�遝Y�uZ/��5��-�˾�1j�LW���M���ݯT"���"{�EB���V`[�37��R'��E��w��c;�뻱~Z�b��.#k��x��}
cw��
����d��j��K(
#׀�e�X�ȱ�c�
s�}���g(D���e,>N��C4N�m��1�nÄ�ryjNc�16��Ԡz��B���~�>��cΆ!��4�ö�[���I?֡���F�$��k#:��צ�u�����6�?��rB,���f�W(���u{?�J�)�F��!��u�Y����P�iP&�6
��O�I��@L�En>��y�k�F��|r���K�1Ic����;�OM1�<V�˿�0�`��	�����^tńb>�[�r'{a�]���}D�$���xfwyy2%9�|�����^�����*؛����g�Z��.ϱV�������b�r���\�d��c����6h��%+�����F1���F����j����?d��*�9Mq�#Է{vj�����'&�g����_���{C`gN��=0���� �U�J�1��A�藢�O_*�X�#���T]�,dbc����W�4]��d�|��sz��p�Qr��R���T��	\K�:o�AI�R�^���7$��}aal� J�mWgo�ݮ�tԴ��e���&Y������J��`\l�g��ܲ��z����p�f�/2����Q	�t�#	y����a-���P!��D�]]P���D�i�|e��I�:B�)�n7����;�&.��0�\9k+U��zg�\����=�)�	�97������|���%�����[��HwN0��`��Yo�$"x+��^}�d��~��A���["�8��^"�n�`�cRx�nTC�x�%TxG��SPī]I�nF�no�h�L�s�����Mkbn� �s���&������9���]�l��
C�� ��l����(�8��$��G]v/�	0��}*�\L�|��'%��o6%P��?/��-�~�AB�4��8�,PI0Q�<�g�Sx��0���Pq��M���RrĦq�-�l9cY�Q;z��'��������vຏϨ�!T���᷸Þ�����`3 �*$(Ir�]H�d��p����emm����@��;L��Ɣ�*�#
h��x��Χ��W++ҝ��p���a�N� WAY*���os�bM.-ҿ��'�g=��]d�e�9g���~y}D� ��+���7�S��n|б�P��6�"$�	����Y%Rg{������k�@̨��O��Lnx���m��AQ���ֱq������!�x�ɅZɞ�G$����oo`P�&�7�W�U}W��D�&�ўL�� �;�#�z2+�O���]SbW@��'�Sb�Մ�H�A�ª���j��j�%��^@
�6�H� ��"�ٶ�.�k4�;�/���?6HmE�4Hq�s~h�.��Zs̡�T<�[��
�,!��Wḛt�ڇ��n*J�B#��kEW͊)up'�0}�Ꮻ��`Q��3 ���;�Sf�!�k��Q�)+H6�{h&����i��JX��3�:M�I'޸�#7��ȏ��C��>Zz&B�\4H�UW_cK0G���.B�~;�@�������+0ƍ�<���9�P���?�AO�SZ�V��h���&�də��iK"�я�QM�����.���or�1m�;ARW�X�cENt��+2bW��p� �U?B�P�e���B��(���>���9Z������(L�!�
?mM�<�_�HI�D��'y��C��o���<|<�T���W^~f�l���	Q
p�wڂ�M����ԙA�Ʃ0"�.�Fet�Wk���g�_FM��(����'�������b4�D��b/c2�Ki�����E�<��uܐv�$�E!U8�����o	��G:8�X{��o|2�f:����M��+t�?:�*QW8me�Oe$DO%���-�mnZ���W����R�D���||��S:����6�J]h��} ۔�ZV U�}7����{�F��A�l�3�FˍD���y��H�����Q����`�?�x'�����"՛z
�s���$���w7�c�%�EL��R��s۔uc���A԰Z�<�+�*79Q�&Lˤ*sD6�a�-�`s�ymsO�jNY�|U����cF�i���a�)�{�.����@z�9w'$q$rpV�f5�:Ɯ��|�1d�9���
��M��ќv��\>:oK�E�Ž�n#�p���Z�����IK��@�`XE�5� W'`KU3�#vj�J=���|�cA�+K��*X�~%�ۇ����1���`��'�L��{)^�k�@�f	��R��oC�X��������8^�v�i^�Å�$�FI4�&-r�OO�J������S��%�c ΋��0�$�`�aR���5�>�}�lK�;���Ǡ}��Lz����9V�tL8�Q?�G����)��Y��
�I_2��~�@���j)�|+����K�f���#"�,�>3̓f��cy��v�k��q[��7!�ԛz�'EQ��Uh8������'�v<~����)v�m 8�^
�l̊�ϓ��-]����J�[S���H̠�1T�ҿ����d9�/�_�]ʑuO�]sAU(a{E����������L��'y���>Af����u�B�.\r�s���'G|*׎������3� zG�uZ[L7t���8�鷴�ǿr˂�2t@	�K
�ۻǪ 0��!��hcP�*�֐������ޥ���ꀲkrTMTz��eN�+�
{-	�zh����`�z��.�6sh�/aQQ�5vVf�(�-8����9�(��L�Dy�.$j��l��Zgb�0�?����.����0��Sd6*������%7�n��"�ݹ=�D��A�bh0�ۯf�˻�d��Y��)�ka<*�+� �	�H��~pu��J��M ���I�EEVG!=��I��p���,�����2�0�͕4 �	
36=7�ho�E?7L�g��p�_�N]?q ��v ��k�a���euP�b�;�9&�QaQhxg��ʯ��6kv%̥K��Ñ���P8��o�騑	*"<���H�֕)����Y}�ɮѬ���m1�A0�p���!�˾P��2*�clY7�F��on�+/�o���a�I�<;P�XŋTZ�'��TWZu�Y^T��a��a��^��@EP��M��KzrEo���m�h�E�H�i��Z@%
��� %��:[yڍj�zh���b>"�U��d`���8е��(���|��'�z�d����kv�=й�	��=8�Ύ��̄�uY�B\�G����3��3�<os�'�<E�3�ػz�b�5n�P����P?!��N|_�?-�(en�l�"�SF�)�Qr���n��uaeԒ�	H���;O�\T�� |�o��蒐���q�o�e6#l:��gf�˴$K��*F��9�|v�[F��V�� i3��S`W����Q{;�^��5�x��	G�ב%���ַL�S�c���w�?��\zQ���tOX�\qs�^�"eZ�[b?�z��*�0�冈Ŭ��l�'q�AV|���5�����~��h�L���0�d��6���A�8"i�)�4���Eل������˭6x�l���˩�NPKe�h�R�Ʈ&Lpei�wB��ṃi�ܿ�qot	
�.����- ��sϮ��Ό�>�����r�����ݹv��刾{��t!dܵ�L���Ge�ِ�4d�h�_����8;�mOc)��e;6�D!���H���`�A��%� ��y�wτr�˷�T�B����>{#E���X����ns�O��ҹ�Mؾ�xЗ�a)�|��6S�R��#A/����)�0 +��"��ڷ	�K�竞�Df�Hj�#�&X���%�o��
_x�ڛ���̝-�T��_1AN\A���,KA.�0���6�����U�+}h���E,O=1��Яe�E�P�:��[�d��|SIN��hUH��b]�j�E
~��2� �X#N�9��QН�<�|
0�z.}�h�&�8���>�{�8q��� �'��L��"JK~���Vi�j�7�V�6�^�tu땩�\{����]��y�F>%d2*P�h�\����R�r�vT~RA�C��CJ uPJ�)�`���=�wW�_C�P��"��ҁ@��(���I
�tK�,Y�gRՃ�c���Q�U��XRA��iI&r��Ep���pBiA:�|v~x7^k�-���Qe��lZ�ޕћ��`�9�ef)��U��F������*2�ޏxH�.��KîM7��"w ,A����+}&�f-t�/���o{,ʳ~_����2�m���Zo�׼l,�%R���P���m�����,�{ٚ��f��\պ0���$X��Z��T��V���@����؎0����f�e���]9����Y	jj�I�Y�w�{`�e��/�ʍ����k
�J�s��K�O�(ö b�`��e�/5!�l����,	�*:uka��F�ɜ]P%�$k��=/X>y.��Ä�xa���XݾG~�l�S#�˭�����[�|a�ZQ ��T��l{~[�]D�H��� "Q.D�*�Ma�J�L<(�LnV+�,����ˌ����5 �J��b�|Z� ��&���섋���i���tj�?���͉9�֝���.�=��O
Ͼn �uV�[s��Vջ��"S���o�^F�[�G��`,�|�D4��h����]�h�@�� �[�[��*N}�G�zT�"����V���[������鮻��Rҕ iy�0��J��WH��޿��Z�[ڈ�9�Gd��=�Q�� Ԋ���O�[BZXAC#�z�~��E}��&����5���nK�����ia���� ���?	��Md���� y�,U��U5<+��1���]`�)���GG�Y�}��g��|�������4�1�Sm~��մ���JE)|�Zt^F�t�&���V����M%	~���^������$}��=���<��-ӟ���F&dc��
l9�͈�T]�ua��Xiw�Tmb�,�O�p5Ѕ�n��-�rzA¶fO�8C�r�}��F ����X68!;���z�hP�Lxs�i2��;B )��� ��\��0��P� �Xh�W���r�ǂ�7n��ς��D)l��3�#�X)6	�r{5w�}�I=��G0�7�"�g&bS��s��R`eh�/�U_�][k�h>���	����l����q�x���J/�|6�x��aq�����ǋ�IQ�V$�pj8Ac���{�tR���8;���H��t�P�%���!��pl)R(;ڽk�@,��Ί�O�3A�	���J��Lb��6Y��Cm��p���Ğ�!r�Ɇ��g8�K�"f�ZV9c��s����	��R��ܱ�		��JU�����Y`��,$��F��I�������rݮ,Ǭ!3��m�iM[W}���h���p���M�ze�F�F�m�
i��*��{�yH�?I1V�p{E� K]��В}��l y��1]�F="T�.N*@׼5p��������㮿bLEʲ��<� �6b��>�tb��.[�������W���2�|Y����Y��]66���$��#�h�������=��w0/'LHq��9B|�K+d��%�	�KfO�C#x?c0b���>$�b�R�| �|�9١3��U�Ů�R:4uz^"HT��l���QJ�.�,{�CP�j�2_�؏Ab��#_�i�g
���j����5���0��L����j���>ݡ��5mp�gb��J��^o�fW3��N���j�'a*�k%�����4��SG�p9��
Լ����u��%7�G�B�����dv�6�v�NR�͢�:X)�lv�*P���M=�&F�c}�A�.sJ�̌���E����!��r��=��8g��rM��,�x��)�b���?�m�&�@1J~�^>뇑pUm�~r5�X't>�!�R��];B�F����֪�V�����W�3&n�$dj�Pv�;���L�8�/R�:�o�uk�+��W �y�9ER�C��s�E������.[+�"��4E6U�,��8�r��'�����+83��Q��B͗Δ��y4�*��������YU�wB�]�̀ker���H�þ��V�&��3���N�_��8L��9���*Y����!��]�GL�Ƌ��>$U�BN����B39Oa4v�˛��<���!��������[@Q�BJ�K�$$} �NT��"�?zv-پ��8�]�!�o]E	����^ǌ�`�l���b��wnx-�_r���:d��,L�m�v��fu	��Vn����"㾨�G$3����z�I���"���쳂V��񕹳�HcpsC�O�ärp�%t�K�ta�*)�i.�F�hE+E��ː��8)"�V�����w�^�̰�fγ[E�z���}\!�%���!A�U��;�v��Eޟ?�����'"4q��x��{kY=��E�B3��h�w��Jߚ�g��uS��`�	(��w���i�g͢�Iu��|8�B��(�s���3[��2��	��.*��R�2P���ǜA��J��)s�\ؓ��eXQ�z��&�` (�ͷ0�sT�K�O�V�����}���HC�AP%�"M��?*2���z��� n��B�~��2"|}�A��ҙ˵;�G�.���
R�Nxzo���;�ȹ��pρ=��P���f��i3�o����C{�st3�k�#KFl������.�����ȳxpiB� ���1`_�Q '[n��l��]��ZS:���bΝչ��d:{����E�]�P�Ѫ)~��Z�q
A5X�C4b�lP��$��b}T�����r!�b�KţB��� ��[?���[���e��Ue3[���l���۵����]9����7�ej�*��:���#B@k�y^q�D�Z�9M�U&�q-����H܆�b�.:	�{�8<y���g)P���D��߉JģFb�i��� �U��u82e�6�M
�b?�9~���M̻��+���h�DPTdN҅[��\�D�ӑ�o�Ho��f��i�A�J�{������Ӛz]�= =��FBT���yN[}.9X��/��c�A���KYrt���T /���P�-�[APε���Y[?�g
�s��V����-S邞��[a�e�����mHѸ��kB�����w_��w��<�*Y�A���\��<�9s�Ajkj�	4'x_-��V��j���0�Y�;P��5q��2Z���,\܀;�[��.��]�<��VD�\�>��xa�W=7��L�6��CG����;9��w�z�vc� ��: ���}��b�ed��"��>�^dsޅaZ\>�ΉĔFN3����	ي��� �^H]!,����\Ze�`����&����bNKN܂�x��Z���zT�q���
��k� ��nE�|�!��37�$/\���w���3O��Q'.WHbn�d���e�9��1�����/����4{9�tMS1:�O3O㏖ˈ<0!�~�C�ܬ|�}�p�|�Px��͸uу�X,Am
ܵTdC��1������5�)Rv[y���a�L~ꈿ��R|u	�U���tQ��*�j��Z�	��?*�� �����/�3��b���o���������L�q��|(��.�H�ο�3��BY�\��Ts�:sj;-�!���`�E�ܞ;3���W3 ���C\1���L��_��X�.�n<�3�#��&d�:��@�0٧~u��h�.�z��țd���⪉�� �Q�y���Kv�H�d����R*i\���mB2�߹�L�������t��T�3͂�/ɟ[��@g� 3��x�a�fý+-�9�&ƣ��&{A2����[0�H�:����J6�)n ���}Mҷݺ� F6%r�~���TW�uW��~�t�{�jU�*���w�
te���P�/�	�<J�w������4�@(������R���"]Q+���� :�����zZ,��&3��O\�X��aIGǤ���)����I������ce���� ����U����ue��'<`R:�0Q0����c�[@����Ґ'^���z��g�KS�o�5dq����ߌ�XmЅD����p��5pc�iw*b��b�`���5��u|�L:���c�Y�ٳ�̱��ĩ�J�#^,�by��%�8V�/�-r)'���v�+���2���xZ|�A�Zv�0[w�VK��2IA�ۆ1vE�P�+n�a'Q��J��u�>��<))�B��"	bF��-���BJw괼\l($�<���Z"�����6�h;!f'�k`Rl��5������u�p���dЊ%
X է�f���>��b!�?�(�L�K[%��Π��2����#\�Ľ�2�/�-"ar�%~n�D3q�D0J��#���Rc[r���=f�������s�����\<��L�����b���ʹ��c���ۮ$g^���YY��5d9#�?����H'�bs�T8	ЕQދQ�CJ���
�h��M^)�����m�9K|sJ3勆qN���O��f$�� U
{P��Hi�v�V�٨Ev�b�ݐ,�5h{�¢�%��#X�h��[�8��{3q�\�����>�����*[��Ol*^���觾Q���,��F�2h�r�,K�F:����r"�<��1)9�_]X���#U>L���@-��"�w\˜<{���)E�݆#8qNbxOn�����q4D�=n��@%�(���8��shӁz��I�V؏�*�#��~�[_�(ѡQ��Ĵ�����r���%�:v�V�kA�b+���W��\N����<]�"x���%�?�-�;����d�'a��VB^�e!D��H���M!E�o�f��J`6j�>�꠽��g���=�0���A�h���k�ꅅ���УC���,�C?i����� ��4ӣ��/i�2� Z�C4�i��7�/L��z��nquA�Z�Kdo�/�/ ���g|p����O�m�_W�h+�#��b�xj)BLs��~�i�f�`�	;P��ԶI���͓� Xୣ�U����:���q����:$�#��Nr��_�gf+��&h���t5� ����+�dm�>	X�e>2��%�%�>2h���̈)�y�gn�X����w�@1��)Ŋ��&#E���wz�1�q;ts���[��"���D��dp+יms�{�	�9�*$�v�,J��w���0��|��
�Ŧ��*�w�{BoR��م���7S%+^�ӡ'�T!-yIN�P�(;L�M�&��SR��o3��b�2sP^4��|�,L�RQӬ�����BC(5�ހ%��a���|zf_��>#�h�6�>"��̛���SqFx�G#f|��`��])��� b�̸M�};���X�%�2�
�8�	���N��r�A
�5�l�`ws�/�9ʫĤN��b� =Vq���D;��t���C3�d9�y��I��P�dr?�O!�u�l`xv&�a�T��ސG��$R�k��T*��-M��;# $.�Y_Zv�^�p�z�����Q$5�[,�&~����Y�=�o��]��A��f�0+S�[ir�o�sЏ72�-)V��AK'�v>�Re_�
�a��znf��%YR��[��t}S>J���>�Ӵ+�ר�_(� *��֠�v�Y�'����!W	� T"?�#��F,��=?�K9d�P�Ӽ*�z�D�S��{��q��"��[�=�N�ҧ���ү����"T�7uUƩ^�zb.
&���ۉ�٤��/��I"�y�d@��
�Ct*"a�tQД�奻'�"��=��"pS$4C^�ﺴJ~|�����3Kt������=
����r%LΔ]Gaq��������㵝1C9(��#�z�֝�*;���I�� ���`h��*XrK�;C�5�ϻ���z���b(Yl�@X�w#����O.���]Gy�����ߪ6��Yz��L�t9����b�mTo�@OW�j�9#נ���Μ)&rp�!K[z���v����yp#��l��d���R��_-�b������)]��g��5��� �&���C�r�o��6ّ��;��CmO��[T}|+�pF�vO}gAh�hgn�w�[K��z0�w�A���G�����d�h�\��u=����9;Xã�ƒxµ8W㹢��ـ�BZ���3)A�X$����e�'<x�n飐��S`�].o����B0$c����s"Uօ$��o�.֟[u&`��Q.2]�M8����O��G{K*& �Cr.��'�Y�԰^Yֵ����ο��1��fB�_�r��6R!PD\5����:%�k!ޞ0��D:�a	� >����j��z�:Ӏ�u� \�1�m����'vǢ�M�I�����f�"}��T Ǒ)����;�����hɕu E+)������s4���3��I�j�JKǥ��?��*CT6��a<�����Ѱ#J�qtc�9��~��]����;�tzct�� ��i5�|ytD؅�<�(��>s��	\�G��O��:�w;�b��W0��-��	��V�`ZO�ZtS��Պ-iF�U�u$� ��ЛfēNhѽ��r�>�]�ǋ֎��6p�O�+o�ר��[;�Z~�;�i.�% u�x�kIl�ǹz�����0���9�G�M�c�Nb����q��6@�ڿ���Z^�� ����n�_���ǒ
4�k�>��*e3R���	�1����~t�Wj����]B�xV��ǬMR�5��(�4�@:�
p y��..anHqY��o�;M�q�_t��lN?0qKh�V�#߫���}e��7�)���WG�d�N����hV�l�A��/� _�D=��!�!`��6PEA0
4=����]�"�R��.�v�u�԰?�ܓ�\�, Y��$����Bw�� fT�W���׿r6{Pp�?�8���=�f�@�$E�D�F��G��a���{����9/C��e!f��H$Y�EM�>Q�w��H�N]����� =!�򰾝�JW3y@?G\���_����㌪��&X4md>�m^4�D|3�b�m0Bt��Vf�I:G�W�2�����d�t��"�q���vf�G�s%M|z�D�"=#A��6�c.�<�X�Ozv�����c̚,�z�|��!��O*����J̪a!uu�q����(R���P�G< Й_�p �H��[As���4\��3������Z)l��h��[�(-��ڃ���Z' ����B`�M�S,�,ʧH�mp~�`=�FEi�\��J���p]�L�:��g?���������x�\گ�y�5��Ð��Ë6��{���w3jy7���K��Iy u�A�B��������C�9����9<�dd>�+�"�'���ғ'$<�"O��G(I�u=��$�Um��g������5��w'��֎��I�Ne��t��K� �$���N��{qFL�y�Gc_���4~b?��n<���A�TFRڦ��&%�BxeS R)�mNh ��M ^�4���\?G@.i1K6�0�q��؎��QC�����4'}�}�E��Z��lr�� �}�r[]�D	IX�V�I,�����!=��od��޲��@�2�^n�q[�\.� �x�m�v�fL�=���®��°�#XhJ�hi�D�%�*Ը��@G���Rz����g���2BQ��#u��I21�Z��:5��}}ze���UǓ���-<�˕�����S��W�J���:���ʂ�?h�Erb�c�	Ң�l��T�e��r�}͋V�p�(Ċrr#�uO<_}�YA7m��Q����%�:�ٗ�0�[(�Jc�NzL�Ls��KADjA%J��Z���m8������8��������yw��I�� ��XZ~�����朅�(����B=�V���S01������	^.)@���s��u���U�LDˀ���?d8���hb
�S�n����"��=&y@��q�F���{�6�g��n��ÏL�3�m��9GήR
�`�>+�x����+�BV������xz���hx3\.gp��Xa�����W�ee���CQ����-jx�4�j�A��"�9��	ܝ$L�(��3T��YϹ����L�<>x�m�U���N ��^��4�T�Ui������xt��a�`�ؘ/4c�Z�J- xA���Ո>J�T���l��?���Q5@��;t�_��ߍ|[tݣ(���+�@���aV�����J������8Y�ۨ�A?[�<:��G�g��ٵ���� ��� ��V	Cx#�I�Τ7� QśC�e������ls�Y�۱������5�1^ W�#��w_��I$V�Nh�ł����pm�	@X��^�Ѓ�moP�)E�qW���$?�^v���IC��j·����B�`Y�(pA��p��"�k����]@iF�AM'MU#�#׽���
��l~~�������]���L8ʹ�c�z�8ء<���[��>c�Uci��U"^~"re�a2�����3K�� �/��#
Qqn��H���n~��Br���-��զ��9��X�ѕLq�)>��MۡZ�!�����i\������`�b�^���:�$w��Yd�\pf��u�_��l�����S(��&�M0�Q����ȵF���8�c���f��XY��&�7������.I���Y%�7].����#�CD ���M��m�G���b�	��Բ`�U����
�3�ř����V�*R���A$& ��Ő��U�C2�..r�.�#��yE�2�'����}ö���9�R�����9R�E	ŐiϹ�wiLB��ß	\զ ��!�h/Qu�1���c7�לC�����H�@;��S�p�[E���N�E�+� 7�uy�)������\�6�0J�m�R3���#9½�~�1��}�i*��ek�NIW�t�?���Їbr����$�����b�i����������1B��e�dH���π-�o,HM&�UJ��3�����M�� 4�FQ�S�f��_��4vGɰ�"Pd�E|˿,����@s���o��ȳf}7�N>I�̻̈́<��P7�0=Vi�g�+,.�m8������8�#x����dv�g���̀�i�H�7SD��{�p��J�T��c�|�?�+��L�n?�"6G{/�������Q����T�0��Ͱt�_�v��z�ʓ���C�e��G!Qc�_��UK��QQ��yT�u�`�{gR�S9O�6�v��k����:ƪ�^�p�fb�b�AR��j%��lݳ���i��!�[�>��a
=���P�*T���e|����¬��&ʦ
�	��;��3q�%�'���:�����9{�H��]:�!��`��N r��h���#�H��k@iDh9B����l�ɔ�H�}6^�i������Ms�J`����s�K�w��U�q�؋��T�C�BŮ5�C?w���@�2���#�L�2��.��CL*v������BU�i�:N"ի5ޣZ �)���D�蜳.���
�Q�_*9���@�m3��C��3Ңn�U!Jdl�����A�p�uɅ}ږ��{v�Wx��J�[�����js��A68|F�h3������u����(��-�z����r�e!�D������J����s�I��"tŏY�(�8%�M�����!���cRϪ�5�W��:	�׃��7o�˹�?��^�<a��O��d���'`��A�̾�Uvʝ��/_q�5�ݪ"T�Yw'B+O�\j[ӯ���S���3q��M���b�%�mod氱�c�Bd($Kj�t_8f4ږ�E��a�2�`��G���(�!�Q �r��ϲ%d�A����H���z\D��q$O�ü�9G���|��g� U&�� =݋G���?�!��	s��h#`�SWd^��~�4�2�~��bf��e�RP?M����46�L	��bx�!��~aI��n%�I�P� t�(vr�t���<\m<��@��uK5zx�T��u������\�˃�X�r��������`ϯ�J�k]�<&������(���!{'.��d�_����#�St���
&m��$F�覺 h<=n)�譭 K�a��G�#G��^{F" >�%�+�Zi�T����KWJ���?O�g�"I�����,���.2xU��B&�D<�m>o�w7rd����dL�v~�!��ߗG8�����%88+������e4�������+�g��9�3ĩc��p^�k��/f�M��6hꈫO��g\��}k�������VG���L���L:�T�>^�M�����;6B⛕��PF�~��v�r���`lp\�@�K��/���P5�=)�E�E�?�@����d�|��H��4�
�/�sQ�h�z�$ha�n�X��-v%4������u
N��=�����NS;	��pi=��f���&�n�"8o���=|�����>��ۋlYy�,�Ϧ�V�> vM����J�pV�h�����9ka\��=��w�k���� ��\�#w���HFS�%!�� �w�	�;E���m.w�i��Pr" @6�b�I�g'fީH^O�CX��ȼ򳹲���c��T7uB�]�spF�t�#�|���3݄U@o&Y(�߉y���	Y�HI�H{{7O�N6K�=Qǝ�&x��y �\��ְd<��w��=>g�o�J}���`^j>�+7��L+�xXRk�/��=�� ��-��fv)��.�Gz�L��x��b�&j����r����=>*s}R;<V}�K#�A"�>:j4D_��7�9��S*J��,6��p��/�>/�2�,7��<3ۑ��X��X�{�(����UG j?F���6�:2f��QE�Ψ/y����>9�+GƔVDz8A�k~��Sٷ&��e�N���L�d�4<�[�JӖ��_#��`��:4�*Xǫ1�p������,s�)F���rY���`+��/.>�yO9|��8fhŠ�;��K�o ��eHt���.2��^��>t�F!_Pn����x]�Bm��T�7��?U����N��a=t�v<�R�̓�hŉ9��>�d�� ����wP$���5�=+� Xm`'���(h��n�gbn5�=���VoS���]�Ҧ�Tٚ�c��6,ɜ$ַQYi��^Z\ӂ�K;��Z�iuEDֈt�aERoz��o�d�U�V�� X�d�2��������>��ܣ�)����L��@oxK��ׁELPBVhoہY�A?p�����C,x��5��cr��$��v�F�9��yTW4v��z�Eݘ���=�T�1���6��e|�f�%k�"#n���mc���8m	\��d��8�]&������0����c�@w�ʗ�}���%� v�I��i��y�7̈́�#��`�\�u�O��f/��>h}���1���a���Z�#�΋{y	��x�Ѡ�����/��x�R��o���܈��tV1���P�����Vc�{3ۗ��i�P�&u��E�t���8���[5
+�����-�j������n�m&��-�4��U@�E��DP�̘�l4�/EJ�D�.�t��v$g���О!��h��,%�{�{0ǨN��C��ŕk����Kr97�_�-���yJӔb��m���:�w��w��{��n�0̴��T�'5�ߞ#/DK�M��6t�G����7���4: H�HA61���r+M��$�H���\u�}��$Voɖ�ǅs
g�ަ�bݏ�� �:>��'��z@-9=���5��J�����$�l�C�3rz������.���
�ك�Y�6�,����I�[�.��~�9��� H{K ������H�!Y�j���8��5pW��1��K�\|�Y��6Y��w����_$
[���!t�k����Q��{� ��7 	_�n��,ñ5v}��F)�(o����3�UA�<��2C��v�V~?l�Tz�k_L`b"��KG�-;m6�P���[�[wR�8�r�riLXG�~fp�%�EP�c�g����^���c`�i!��h��y�ҋ���r�G�[u�Ē|OT�h0��k��Fܕp��Zj�齢���N��X�z'4İ���){�ǘy�#��~m��y�,��ڬ�)�����a���$�R��e�"��((n��|�ỗ�1}X�!)!E��j+i���Ώ�!�����8Fi��~~����kn�d�81h�m?����3ĸ��'�+F�y�:�������� �Gi���%��~i�F�R�W��ٿ����
�K?�8�XmA�L�ʅ����b�8���sG8�m�4ڪ��j��v���r!�t�4�3����rx� �/e��a(	r(k��X�M���C|�L�;�}(�@f&W�y��an���X2֘rtsYmk*5P�y6�CX�mߌV�<�����(���e�vZK,�v�/�ԧ��hUD��3����~�G\�j�<�xpxe��JLo��B�#�
��:q��Y�i��6K\�4~�P9��.c���J7�����(Ǧ�f_�������$�]�z6q�.ǐ�i��#�50��{�JK\S��Kl�ރ�^l��d!Mt�s��nh,�N������r��J���I*���U�X#�oă1��2:�lo��ʞ.�Ǣ [8��j�=�����A����`٥A!rp�!�U�x��8���R���ȅ��Koq�z4[:�)�|��{J�i���w�]"N=����nC_����M'xS�4?�g�=q*(�齱j>�+ׯ�f��P���������!��߹�K!���dq��l���q��,�=�	Lm������j�V�G�����>074f!����I��W����|-(&����JN��D �� �7' ן�B��G����a�����RL��Gk���-c���P�|�_c6�~���F����i��<��d/�k	��k�KW��Z�^���p���a5x7)�m�V�uU2-�1�,���.����+(l���+����|,��`lIU��X��i����Ʒ�.4���-��0�"P�+�|a2db�{^�U,J�ǓlqT��g���l���Z�[�cͪ2�g�� &D�kPu��������sC��T�>��v'&2��Z��c���y���^v@��r�Y���e#N����p3�F���ϯ�a���}-C���[�a�f�!�NJ\��#��3Rl��_c��Z����7���IB
���0�俗2�-b��	&��I+����+����b����=���bx�6��x��U�K��2��_�/"�Fi�gl�%I�\�IlD��%в�-ũ<]g�3 �|��'>C7��v��*yq�#1zwE��*�h�w����n*,lrxvJ�v��g�_H�膵1�m���;���"���f|m;l�Y�-�4_�	�'<.�� @)��ܝt�I{`�إyȻ��r
�_�C��6&�H�{M=�i�9e�{è��%����Sۛ1���0�� G$��&���!O�M�C/���Ӡ��,B��&���)������<�k�c�e�w֫jT�V�!�Ł�-	"M`�W��Kd�~~��i����6������pD&��"%��P�~$u����
0d��v�1��� ��{��H��C��F
]�`�Ox�orhQf��Z�f�W!���MJ]�u����.l���r��6�4[�0�ug���zS$���A���!w1L��Hc���u��v���K�{�oOe�TGs��8�f�v3�<7x<M��,z�)K7f� »U����5��$K��K'[$i��e�y���<��l��K%8SP)�8W���(Ag@a`�݂3>(@$��P�J�����v�,�X�c��#���B��.RjST��=鳵Zּ�90�uP_��8�>�_���#�z��p�6�L
�ZI��J u�������p�C�9�#�\�_j����OO;_b}�a�,G0ܕ����i�G�dӼ�6�,��Σ���e�8�d0bh�;�)�����Q���ԼG'�]��%+D��UCrŌ\�(��.tr˵���$m�E	rJGiO-�+j��dF��7yS��t��R��?�Z�u�R�}�Af���(�$��_Yu��~��n)�=ۢ�O����޺*�u�gm�y���.)�b?��š��@��h�(�f��#2�r>$�,�aj�{|ХeZ��E�K@�$��*�`�Kx]�+'RN���$5����:17��!��}Wk�J�_@�hy.۶5g��˔�h�6�ZP�lئ�!*��o ~��N�G���+y�
Ժ��}�K�v�ߩ+��Ԯ0|0']���x.+���񳇄b��	��}�VMV��Pcf�����n�_�fC}��4��p���^"�&����C��*f+z{�R�g��آ������G����9�y=�B�ו��톱"��lR%m��J�|���#O�ZN��okyh҂��z�%;5i!_'�%�É�|��J�H<���C7��h�W����ddͺ������J���!�T��0�D�<!�&�'�8�Z��Ww0���$�)� g/<r�0��p�5���`N�_�G��KN��\
)ǁ�;�I�������#:���!� �Ǧ��e�ZZ��}ܿ��zf"X� ��l$�4/���C�lc2G{N��N��^�a�m�j�?�\uA���	�}P(.Y0��<�T(�e#|�����S`~)��i�b���Ĕ7�Hh����a��,҃RY	%�;��.u`�O$I#��p�C��8縘]_e�sͤ�~mT�j���/�FІ�P̨��Y6���U��#�|���<(�,�o� �)�5�[x.m۰���t��1v���aVLt���D?�:Ú�a����5�i�9Rj��sq��o��Ah���v1�d����n"����J���Wz�,��6���#�{�_��(V��(Iѧ�p���s,���mǬ.,@!�4h5�<OsASy��G��A\��VL�-��+`ew������R�8,��ab��
<���Ŝ�K���C�����W-ʧ�br��N+�zf�	x0�$Ew/ZTRq��wΔ��I}B�}׵���e�r����b:�0^Z���� Ⱦ�%�C>��8�5h�bK�����]��/r_��'ɳ�ɝQq:�HI��C�<�<ͷ�3|���oH�X�����,F�룶Y��M��}T5;D�z�(e�:�3�@�(�v5�X�`�U�CO�GN��4�$Av���Eu�`;[ �=�����C�:H�Ì$b���bR�0eI 4ݵqW����/�O�v��9경�]�Xt�xJ�pQ�+0��-wsc�c�E^j3�!� (zC�Gb�B��@�bq�����M���������C�l���~И���|Y^H�W�l���Be���ɪ�RV�J!����۽|?A%s�>�:zOs��^[���CT�v�c ��vJ�l��x���,��`���N��GrU�f����p\��@g����
�ud��#�S{{@�c7q������=�:�93���&���-ԉ;*B�����R�@�@�K��8������a��CO06>�ZC�A��RUО���Wg�ж�{��l�O~��bA&+(n�!)k:�K~b���s`��yjCxP��&�R�U :_�"HF`RI���6
��:-"z� ,g���Xb`����2E:���7���k�In0��Os�S�w�f����D�	_I3�ۺDmܻ���)6V��f[9ŌBP�ΧS=ˬ���X���S�ҍg�@&dn�?�(R9�a׳�|��]9�`��L�M��W�c ���:��Q�`W(▸��'���3�{�¾���3��%�"�<���WO8�y'h�(�}�%Ʊ��9���tS����¢=|M��-G���G�!d�Jш�&P|���$����)��`�{���J:�qA:'�y�~�J6�d4!�a[��x��ɑ�R}�h�y0��&�Zl"̎eU���骞�hil �+��!d�}0H�)��"�>;MfZE&�Қ*o�t�5^:i���w�?��no0�Hp.����N�0;��S<�:7w����T}�������֕�\<l�4ġ�e�_	
	]:�Dv�|� ٮ:��|�N�廑s&�����}��D�
*���m(����jk����אO��ZUd���Ǣ�q?]���	'�֟��4P��L'��t�F��rɋ<ı�S��h��E��O�7���B펾��F{*aez��U!�Ƽ�5�������cHtk�����O;��T����MdyH���*t�j�v�ῑ3��)
�zzz��z���N�Pf�c�Z&���S���Y�Wՙc���:�P-�!��ٜ��!R=�AXp*N�1���t`r�<�<��
���3��ï�~Ǯ̩:�ૡ�C5Nia�x�/��A��PS��3���Ma�DC �|`
��x��(l�;e�=��3b�L�C���]��ޛ�E�'���	lH�r:�`ie� ����P�2|���[����TTqr��M0�Gi^ֵ��ǆ��-ʍzP��e�}EF���F0H���b	r\�4|!�o�|DEmt�s�S w���b�Ͼ�/g�V��.���mo�؀h��/|4�ED�Z0�on�YShd�p�n>�ӱ�K�^j��*/�I�Ն����7��q6��9�p��i�AI����0/��k�|�]��ڹZ�8��|f<�$���Mx�<���[��$G���������b�~
d�B�e�!=�Q�?��^��@�)�ՠF��gLC��8��gO4�g��܏ƻ��cQ���A�\��z��vR�1;;��?)s(�g]�p�����9-���~���*�~���x{�^\=�v,ѩ��_i _�l���|0ljA��Z?7	�\����	���3�.Y�H�Wx+�W��E��I� 6Fn�S��#��(%c����a�<~ײux�	3L�%@�
K�S>������Y���.���	�q͏FR�'q���C4��
;>�8�#�x�xYjO���5Z�9���W	�U#�4}��#��m@	���݌�}8��,@O������G��o��l f �:����o�ܣ9�Ԅ�j
��b&g��ϕΤ��%���� ��;���
s��J��*D��
��U2�8'�y���=B��f;:�����z��ݴ�jM�u��#K�������`*Nec/7��!P�F�}��m��֨��ԺB.ߘ��fm)� �ϽF�����#`[��eg�?p���@���Ϗ0�k�_�U�N�<�nTS����A�O4c�	��-s?�9PWԆ�!��>R�q��^o�k�z�lؗUA�8��6*{�J򟏔!�nF}��z9��'0 ��k��EUS� ;>�18xHJ}Fa�}��YG�.K��`n�|{SOT�'̵���v 0I�,��N��F������X,����(�h�X��o�)Gw�X�/'P���k��)�7��A1~J������G�3�`���Kv��r�09��7J�H�]γ_Ge�z�G�yɞ����8��;���ie!&F殽\WSl7r�G�?�8�9���jB�~[x��Z�ȩF�8����~w¦4�^~bv�m�+W
D(f��L�_���~�|��c�8c��d̍gI����J#�E�K�B,�ҏc��MI��S����K__D�pZ���,FΚxg��p#Q/�b�S������cJu6�;s#<^�����i�|��jVG���~�{�a)����&D�[<�.l��r:�t59o�^�W�q�?���<�d�����pdu ���*�͸qLp�fuo�x.�Q��CdeA���>JP��R	6���J�"�,~��"�[;���o9U��~����}�E,�e�7h.<9��D���*c,�gV3��L/�_h��ޜ��}�rWˊ	>�9v�LNe8	f�?�&k}J~���c�a�a���� �yݿ`yE��mE%|�?<���n����	�dN( �R��Ր��,���O��E&;�6MtW�zJe˛.w�������S��W�^��P.*�g���"�N�\�v�A�W.��<		ӏjH�y��r��!��F�To���������}]�b7��	e�}M�J�� G�b$���|�og</bn�i���D�u����\��X�
�PJ�kx�6P{i��k�*C|7"�|���<�����q�`�Q�U��a��es2�u\w�Jh1����K!����"�P���P`�+܁Kz�s��4�ud������͉����b��z�5&:۔��5�e��,��k�� �:!�6��D�/�J���Xtv�i8��:��z�N
9J�h�w��Z�\�N s�y?��s>�<m�t��x�8�ʜ���AL"�����"��'�t�p��|~S.v���w]U��}SDrY":�5���iK���*�mQH�I��f��o�v�&3D��t��"�C-�O�*�F,✻��l�%�w�8d��B]a���4��X�M���7(Z�" �%,��
���S�>,_�41�c	Ը��<6 \��޷2
<O�j9���>�vZy�n�fs)R�1fm�-�z�E]�4mG�ܧΑm��Q��wO1���_���Њ[��:%9b E�hk��8��exHȤ�I���?A^�Y&�iY�M��U#] ���R�pt�O�Hc���/\���J����W��6L�GM=��)tE�>�j�� ���1D�E*��n��pSؐDԏ��Qh>��u�Z-~f���@/RiF����M�Z���t@LE.0�$��qJbs��8*�İ�_+ik���ͱ���lЬ�vi��1 �qq]u㿟��_�K❓�#' ��m�%�|��!03�E6��F��kr$=��d#f=�C@���g���s�zw)/|��ĵ��گ�+���]Tԣj���5_�R�u�yQ��Ǖ��7���1�evi����J�Y�#��e1B��vQaĨ�2{l��͖L�0�����4$��j�s�׉F���X�r1<�)b~.L8!$ߐ g^4l���웟L'�~��u_b�f������`�f'��fA2jqm�&�q� ���ĺ� �6
G��(�@3��1�x�`g=>$$iғ���0�� dƼB�������lT���K"0HWt���B�s�����2h/���V;�^��10$�l���M�o�(���Ql/��wJ	պd]��۷@�Ρ2H7�Ф���dQsC�t�}���+>%z��l"��kwI/��*�q2�h��ށW�6�1.*O�ΖD��� �;^���^���t�?3�Z�fb�#��H��@�"]�:8f�4���[��&
l�Y��:����_Tb�L?����M�:J�l�GB�O��?������vVKAbip�p����	ԹqAgɬq��n�d�|�
��wE�
��Se�J��,�fa�Z�2��d�U�	 	�U�j�A3X4�m8�yi��px�rj�)��w��m���EҊ�k���WOV��g�$Z�(��R�%迳}�,s`O7�|�ى�co�>� 3�ͧ�^����V�:�	b�ԏp 7t�F�O@��@��7�Ys���=�W8#�V$�-���܆��X�K���?dٔ|�X��$�������M�oJ���:�Us��
�\oSO�.f@�SJGDA�I�t�D�B�H|P�]F�kW��:>\'���.P�;v���Cw����y*D���i��f�]�t���f�]H��Lp�( :�K/I"b���U7��s|d��y]E0�9Լ݆o��$�+)�8u|p�N,2���I��O���Y�gv���7Dnt�\	?[aϚ��]��,d��5[�����T,�j�'�6���������?�zm�3'��)`��s	K�,�Eb#��
0�,+,
���1����y���6�^&�S6�P�Oz7��Si�>�&F�u@�Vv��um�d��!����G������(q��#��oI'���֦�3��r��u���7�h��su2Kp��f��.>XM2F�lLV�n�
�+e��%<��>����(?ٹ��e��)Qէ���7>~��)���I��D�`�BD��_���n�nM�*��4�}Ǌn�At�G0� ��{�i'h�*!b�~?!��"�\�	]U���Y,�rY�=ۤ-N�2������!�x�F��p���O[�N���f�Q���?��s�GkP��K�X���e@��b/2��ďQ�R[q�{�=�M����Nw�#�7�	�>&�8S�$�&�̢�!��vG�q�5]���ƀ���>;���+�'�)����vw>�d�4#�T�,{?$g�r�0�ߠ�\��5)���9��-�W�J�o]�ŅI5Y%�P����j�����s�sf�+"�hez�'��� �$]Чi�& /=��gVc$dׂ�T4�1�t[�O�M%���\�Շ��6+	���E�:i�P[��n�n����1���=���b�x�4�j픩m 3Hgu5$O�wR;v�5V�2�x�٦�Z~��k?{5?zҹ�W�>�7T���P���(��/�^���<��/��vآ]U��~h�q�D�ȝ�,R�x=����Bl�[G�2�,��q&�hQ��D�i�T�^�vA��1��Q�j���\�*9D�|�����;�"tt������QD�־W�����h����1����Ď�S�3׎0��Q���tU@e쁩̲�s.�34t4����ډW�o�}���?��/��?6<볠��g��,���I����b}GJ�>�e��!�
��S~x@7)�~��s8+#�D�Ή�Rp�Y�L��S��&��~g�7�e.����4�2�mT��@�f78ҹY�rW�T����𭣝 TEOK�d �#4�g�챻Z�����Q��}��o��?-�|��f?�X���Z�M�=�woo,a��E��z#!�@���D��B,T"�Z������l���j}���>1�zK�kt` �E~���B�u���ꩯy���WufT���7Y�Z�^��ߞϜ��Z�2�6Nq��(��z<9dpO������_�ٙ�	��zqؿ���+-�>G[1�� &���
r�:�(�SB]d�) �pTB$f|	n����u��J"*$���$�ZA��y����/N7%J@k�E���9�����&,P>*@8M�|Jq���3�E�&����x�5�>��݋�O�j�T���]R�Z8�1��������~��K�sb��+tj�E9쏊���k��!x�c�tC����Zw1��Ʈҙ(���D��"f�^�!ʑKO���@��@��!@v������@�N�xl]', ���Z��!�٪s�����]��d�Q����?�}�3?���B�?E$3Kr���$�<��c��6�^��&Ƞ&��t�Ga*���l�W]��LQ���g`H�ڵ���2���3^=�3.�6u�0�I@2�P5y���A����8BG�ؔ�^���	�dj���f��>Ue�t������U�>��^B��yt��w�t���.���i���6�����b] ����)p_$� ~�ҹ���a���%���WʸS����!���rs�a�v��
�A�z�m�����������������d�nB�����: _V��mn��e�^ʏ��펤�E(u�r�Ý����E�#ߋkz
K���$��9�$k�1���#F�w^�O�f�6�xg���э%�s��7)k���r�_�ge���wӈ�Lݎ=���#�$���C����������U�:Gj<�?\C�h�k�<��$�B�w��H��D�C.XQ���?S��7����b�x�}��[�5B��K8��>Y�����͎��~�շ�N��<pl1�o>RAZ�E���� �@� ����0:�ˬ_�6&�[�O\�B���ѭ������,���9�H`�4�-+s�Hg�COo������"���Ū���Y%�}���V�=MË^�W���3��倄Hm��'�oH$Y��Ölҹ,��y�
)	"���=�٥}C2��נ?1��в�o�G�o�p)�N��1�����/8�{
�v&�=<���{[��8��O�lqK'�i�}��n_Bv��!m�G������Q�Y�2�N���FQ�&op��eWk���(��1"g6��
{2T�|�g�?�ȼ����69zMy4����Í2ǡ�G��!����qb��T�qE�/8w�O�Ф�iK҂F��}. .Q���ܖ���hf�4�������tl�Q��6#�笉��v���ﯞ�)@or'C�;f&�ieM�����_G�eڐ"�AQ�Z%GY�iT�IV���N4V
Q���a,
>ъ��s��G���c�N�L�|�Qc��]��K=-=߈J�J�4�	�
�����h����A\��R��d�{��T���A>�1?���(�ma�����i��	����pC����#����?@�'OU`m�#u�O�^r>�(���*����-��V�9l�	�tA����KM�/�U-6�/�0�j��i�K	Ʌ4	A������;/���ey��D���Q3�:�wؙ��Py�!��G��5�a��`��rk�~�m���$��k8�p���H�"�B�8L\���0�P�d�!��"t�[(�;����â�]�2�C3�Z�3���r�%�a�j9��~r4��3
��`�aY&�y�WQ9c'Q��:X
�;qeS$$$�ڀ��u�/\�[2M�=$,��xH�Թ󅽅6� �9B�����V/�'�P!����A�����x�&���w����s��y�z?SNz�9�&�Ϳ5 �N���<K -t���>��9��y��]�dz�_�=C2���wx|ޭ��M���z�%��&��^�Ղ�b�}��� � �\�9�o�+���&6M;rOm���u�s.q��I����xx�bF��U��50�uD��"s;����%r�Z
�6�]i���O�TL�YMhL��y��n���X�Y�	�Ǚ�#)uP�o�MY��,*�6�b��=&������̺���^&Z���<�[�?@_�:,ix� Ȧ� `W� �}f.Ƭ�����H���#�CN��N'.#SM?���0����#U�����WyE���w#�3��Z�%�h-US{�9�2�[j�Y|�vV�)��=�.GV�̷�KQTS���/����E�{Z� LKloñ�|o�Z��Qϗ�"������D܅G��J�a�DH���Xj謽��f>�A�,��tt�J6'�H���)m�=M��z
k�5�1�-n��v*�] �lR����T0�ܤ���w��nX�v/�ȟ��Υ�SSE�}MS�k������D�WbJ+'���hf��ۋt^���f����k�_]�<A>�q�i����>�{�2_BLv�y%k|ЊOdf��V�Ju��n�liz����/)���ީ����|O*�ch��1yo@�Z�Q`'�q�#�4��d�j��
s(�f���Q��*�
¡�&י�ub(��;�m��d,������}�ii~�~����e5>�-/�2���"��}�B]չky��%Ci��vӄ-��?�^���~w{��&��nJ����i��YnqF�".uB����`��^�8��1A��l�(^�o�%����2���@�� l�ُ�����2ȉ��Wb2[e"��'���8�4r����b�E�K,��돳L���º!K�W��֬f�+�����Z/?��Tk9��z�/c�
_�:d��� 4����l韞�Y�{1��O����o+��v��Ϋ�;��-�H�5�uݱ^���t�R'�LG��c:]ҵ:���g�1�nͬ�,��/s�|S=���3(��~�bH�;�.B����$z֭l� h Xя J��B����������M�]Ԓ�:�Cε���,���r���Zc���LZ\&.�eIIR�+�כ֡+�OQ���ߖk9[��nP����/g�L9�ް���+�B�>�^Yr�����9�x>$?���^��Q����D���n���x�	�c2y�������p��a��7,8P������qԑ�9�6~Md�p
Q���o���u���/���1e���b	$���^�c�"oO��{�|�	�_}Y��u�'XwH?�;��G?��k�>��Ԧ\�	ϫv�o����'\�8��%x�qѸW0/s�!T͟�i�,��'F4��[�}��;V@�J�\�.#�a��`�2K	U�o�8[W��H,E�$\�t���
�:엹W܈��(��K1�(���|L��&/��ߕ8L�;���|Z���!W��2�,��������l��>�l�؋i�ȟ8���"q+>��m��G�d�363 :
1W ���K�}���@Y��<���\Z����Tz���ؖ:v�I,�NPKc�uq''��>�n�o���݇) M/�-�b�]��Z�Z�Y�y�6���Z��#�pX�Rl��8=�ϗ���c�U�+�����:V���)����)��O_�c_{Va�F�x�t`t�)0�x6�� @�W�ifg�����o��{A)#��7��"7��hk��	4agn��Ğ2x�2�c�w��;�綳@���9����Ր���dyiN�}>60
<BRW��QAm����&��%�Н ~{^��}m��%��%�[�H(��Ģ������-�f>�����'�RV��
�ǹ�~yչ���������"ŧʍ��tS�f�˪�w��{������&����;p[���?¡�e� 1?T0��0�$u��,��	L��G�Ut�Mc�.o���2{�:t�XH_�{��
e,Wj��2�!s$ȳ8K[�=/�6!�)+^"<ρrR���˺�mF�m��1S�&��^O���!�M�M�%�j[)ā��>���c&qs�@k����<,dT�wN`f��W��"^'XÎ�*q���}� ��=?:$�_��h��B�ld�IpI`��3@ax���Yɯ<��T���a��6&Xd����_�}���7Y���PY�-[oJ	�|�"Y�j�JE�~?#Xu��� e��oh�`�����Oek/®�	��A^�\9�WAb�.�������\_��0(\3�%3�k��@#ѕ���a� �[��sg�g�w�-�-�|���0n�v�@L|�K\�:����h
���E����#�my!|.�G�{�x}IT��{z)��%�X<)[���_V�&����	罖-+9�j	��Ȍ�1�7Kh�"ť$0�����M�Or����l�=ju��֖�S�-�������^�,f�H?K��p��^�34Y��΋^ͺn�޽�oLC�v:�'�}[��:n��������)�?D��<E�&�[tZd@�d�
�nѰ�������|2Y�n�����)���d�猗��S��ܲ�SI��z>{���/�2l�^�y�P`�a�y9�RIA�������u<��T�?_ۋ&�m	A�֥�2�;�/�H��#��k3jE�_M7G{)FmT�ꋖՀ��-?����/�ֱǉ��/��W��v�̺e���*��F6��IE��W/S�Od|��Km��8�w3�"d��Gn����IQ�DF=�	Ŷ��=ϊ�E������L���Z�V�"�C����[��wM$�j?y�Ti#��hs�=n�M�Z�q�tLO\ZH9�5�qW�r��XM��!�^Y ������y�<�ߖ���k�(�a��r�B�h@R>��1;���
�k�C_5J�0"��0jh�����X����\9g�ע�z��k:	�*�2M\Pt�~�E��f��O�iIH0�[Ӕ�9�*�˔U��/���>�k$L�*D<T
�������@9�Y>k^L4f��m׶DS��h�RS$�:�/L�i!������b<[�Ɠvv�:ǤɋZ��)SG��5w���4��i\�.#�[��̖����`�5�����H�?~g#�Am�
Y�Q6}.H���5�~{�:ȸ���َ��e׵tf���C��I
]��c^A%���ϰ��L���ܰ1�z�1���j6��|E����L:u��J�=����N�((F���	^w���:����l���	�}A��h�2��.#���&M�O�d���&_B;o��I�0}����(�� 0�a���d
8j.ӯ���c�i���L3K�H�F�c�����y?E<��dUZpP��������4!��Y��h�y}���|�Z�����0�G��}�}a�����N?�t����'O��xjq<�8���N5�V���&�=z��}���c���)�zw��S
jt���$O�g��rвѻW������tɁ�dl�ih|a�W¿/n,� ��ퟗ��0�m&����Zgn�0]�?os2R�]"���'�4W\PVz�_l�"a�G8���X/�����r )�MR{I��Ln�<��T�'_�'��L��=OC��Y[M A}��_����㥺��
ջ�m���W�4�;%L`R}]#U]��l�A)UN�4���2�Nc��� �Z�a��I�yj�����:!Y.��7v�'���ǟ�*�t����M����^+d��:N���^4�RuT���B3�s^3�D=#������4��NR�S� ��	R���m�_�����d�{��4��&O|mO{x��@��qXQƠg@�`F��\�PE>Qϊ4��{<�2������UW7��|\�t�S!� ��3�
kɆ�2�h�i�:��!nc���JBC���!��'�,����/R���,1���Uf���	3C�䲿�<[���ΐ)B��NcS�pu��{��dt��%@�7
.�((����#�C'��S�h��Ls:#���70��ēPr��Z����3�qCQ�BnѾ��+:���@nQ�p�<"t�S�"Jo�6�NJ!�WX���/0g�獒�A��C
f�<c�@N_���/�f��BGق,��מ<��P޽�qaa]��*_F|�c�afFD���\L�/�h�C��V�2�-9����(A�`�������[~�2FБ��ײw|9�7���*љ5z�y���\(�u۽a�rE�/j��Fv�p� 1)7���I��-�>L�L��P���a8�R|�-T]�;p�`��- �&�c��M���uݨ'$�)��j�U�-������,-��4�vނ�jO
[�I�T0h<�B� �4Ŀ8+Gr���ewo�����/L"'Z�Y�Z(h,��Š�y��c�X� �u���
�I��w���R�5�R3����6_E_-#Z'��(�����1ȩ
��ꍸǎ�0�b]�o!=������U�;�鳑��_�o\�G���#���a������h����w����+㰿�!����c�����M��or�@0�A�"V���ꛋ�o�|k�~�q�T�"U�>�u�4��)K报�}��]L�zT�w��$x	]-Ԭ��������"��b�)�oy������+(0��%�����I�x�<�~�&-�^M�'��~Y�{��iX`p�}^�_5����<�=B�֔�t��8v����\�< ��ECJu�chk��<��h�I=PUǀl�/��u&�)d4��r���Z��*�N�1-_��i�%�v���~����륩�<����Fr�*�<��ݺ�;�(ٲ *X8Tm��j�i�6Ԅ�4�Q�"��輣��A[����P��ш*Ж�BTi���F.g0r���I�_}(+*~�j1|]��ܨ؃��fr&%�I���Ap��[��Zw4Ge����s�·�5n�Q��F�ӥS��ny��?����7B*�r,;�j�,��=M�X�BR�����,t��D=`�mv6�m������q��+��}�"j�CY��v"�l�➂~8/�#���5�B�9�;2�jS'/�q�D"x~ܪDȚ%&����
L���zt���+u����m`��7��gJ�V܊�5AA��]ӷﾮ�{��9]>CO[���`ܕw�����D^6��@�$������p�'yt#W�����{M��,�֥p���}N|T�0��Y+�����n�_m�
�J�=�s���hj�	q޴4/�������H	��x<�?��T{|Ѽ^�H�+�k����[S/��$mb�}p���-8:�Pt|��Ъ�����w6�K��v������y��-��"�����(��o�� �������A�J�7� E�cb���R6� �"��+�󉥄Yrb�(x�&���x���������^:a1՝�ƹ�Z��n�ZK?�D���w�F-��O��N����bC����/i,�]5[��O�p9$�6��I���LK|��i���4�0x@Û��h��P(�E�����i�4dX���X�\�^֊s�`-�u$��f�->��lݛ�����R[��^�wڌj��8�x	G�8�H�2���!˱� x�`Q����5@Vp�Y���#ǂ�z8����O�+��!�R�9�a~<y����k�L��� �s�8��3j�MA�-P��-Z!}���"�2X�M9�B�/�Wmw`_Z��Fe����4H���x,�W�9���2���Լ"�#J��t��R�T��5�{$�����PԶ�M���������*�x�����A/�"瓟�7�u��������"��Vχ�v�$��s�����"��z�K�k�->ӧ4�bܢ�?ɔ���;���h˼�q��:�D���IQ϶���ܸ��AR��P1�Lewi�����=h����FϪ��_1&��l�ϯŐ5O���'�T�� K� +��φ�������Y���H7�z^/&�sk�zɂ�^J%�c9QvJ�i~Jy��4�`��8�#���������n���!c߲�{;��f�\���М�^_pg�sw���oɎ��d�a&$�^��L'Ѡ�C�τ1 �D�v����ۡ�a�d��Vl���z��"iZp� r$Ƙcq��M�:����������'��`h���Z�~+�?��ȕ��K]	.jo� TA�d�ay������-�0��4{���L{��~�H{�c�<�9a�y�ן+�V��b�Tx~�/����'J�-��A�r�{4��Y��'G	���q4�->a�&\-q��?�W��QF~s��q�t>2�;��H,�6���%6��N>���u����i��k��Y0�"K��%أ0h�m���ѝ�Hzǘ�h�AZ�[Y8�eC
��
J�3�(~� �ZoP����)�u5\6�7e�']�\�������6��I-��ɋ����D~ �9U�G��zQU�[�Sί��H/�v��-��o�9D��(ʱ�� hQ�*����V �qE=g���ȳ����1�O�Aݱ�k0y���,'!�5xV��Bu�<m�f,�{�`�w.�|A��0������N����g���y_�������|��Ƒl��s�<�'f�_%Vف�b��:��xN��0Mn��y�Ij��|�w˄*�vo�^�,v�c'�n$�U �w[�90��S[Aq�~3�$�~�Y��� :�f5�Y�=�Y��fV����o7�&�,S��M �T��p�qщ��jn�Rz%ȔCm�5_��z�~V��%:�п)�y�@��2�� i�G��p)6�
��k�NP�u�+`R����+u���O~�C�R�%udl�ua�%U����i�D�T��lvrA5��.~С���?h���_w]á�`�1����s����0��/�Ƞ.�kf�[�C�͆j�޲��V�G���z $��X���~�gJ�<�Ȣ��u�ěo\��3�^1ˤ+2�/�J���hV�&���F,P�ZmoO��*%�}�X�Z!D����� :�z�Z�d��k���W����I�v�v��L�ֻ�yzH�g�euS>�d�@�P�	�*A�D@.R�	�Nic>���l�WC�D(��<�6vF�+yw��C:?}y�k2���uY�(c��%kJ��#�m�&	a-��HV�*$�q�!jffyR����X�(x���\�K��gU8�w����[�$�Fp��W�טJ�Γg\ ���R�Hzz^۾x2�i�NG"�>-�i��;�Bֽ�Ơ�c",�{Kd������.��r/Ec���x����&]�W��	�f��!Q�}R?S�C�#.��%����0-������Ľ%.�@������&���Q��'���Wk8�>@)Dm��u���fD�.�q��"�`9-��h�E��) ��S4����망����|�P�3���d���w.c�8�@ꊕǒ�)$�n��������kV�
���x��hj9�A��/�1Pu]��^hc����Q�Es\�L�D"<���d�'&�.3��-[P?B��&�{o��LR�I�r[p�Ц#p��:�$���?���9�:�z�7��q2�ɰ7D?
�'�~\I��*&�O����fx7<d2�����W�o��"�� ���T;\QӁ��	��q���w��x�!��nɀ:��h�
B�@Zv޿$�����.T5�N���gՅZ6�/��z��5���i`0�ޭc��!�u"ɯ���>|!"kO��6O�9F���2�}{z��s�m��wJ3�
�Q;���獮�9��%"��,?�]kVAǦ��
1;#W��&���i5�n6;6j?�G�Srg!�tGk�����R,1l9V �$���4�,q��cۏr��P�ާqp��W'_*�1g��2�e�f�.�rmuQ�ۚ��wj�᭵R�c�BFu*%���Γ~�X���v�z��yn�S�ڠ���,��Z�`��-j:z�-����))LF>kW��%H���}v��#]5��7����Q���d���-���o�"�i��E#�u�}�8�D7�Gߤ<���? m����kJ����!��Z#��%���0gE�K]R@��`ߢ���x� C���?��/�Kc^��i�VJ �,��=�k-�]�M�=��C���q]<6��k�2�_�)���7�����R#�\(����X$���[	���o[g�K����-�!4�E&r��q�����\ܡe:�#O��/���
SPvDSx�
���|�ק�c,�f��n��@�Y�{�����P���zM�i�Y�58��t.Bc�����$��AW�߽ޏ�!G��:��洞�a�;����Ag�%$���DT.��s��鄰�����LL`֔����O"�L9��L�K61��0��<&�BiDt�簶=62��]�F�-_$]^�����tL�?\ߑ][�ӓ��ࢵ1�w�����fǠQ5�z�C��уe} �� �����sm���P�(2i���R��L��6�s	����� �]C�~4ӎ5}�ߓHW� ��sZzZ9��ƅ^�Nf���:5ˇd��G4)B8�qc��+����ǹ�Sʧ�NB���n��� �2p
�ABc/��H�ah�/p��j�!���
Z�z�V�i!l۹f$8Í����E�m���O�!���7��U�$3HIX�bt�f���*f~�mA�`�?AT �P�@��¦���S_��2�?5��x��WB��^��g<���P,�Q������ٛ� }�(g�K�r�+����&'�_�Q<���@�&�4'��wcaF�!nC����lt�>��#.nֵ���+����z1�& +2X��h�Q�gd�*�I����s���G�����l����a��؛�T��)��x��1�L��R
D.�Y��衠PXQW����	�p��ղ`yR�P���%�x��hv��G3�s��2l�0E����r�&���Z	ӫ᠀�қ�7�c	�Ɋ)93��%:�K�Pg�Ls�<Eq�M2d��W]<;F
�j3P��E��g�6oADG;�R��QCG��ډ_d#��g�(ŋ��AI��*)��Ct^�Ng�{Q�CRr¯��+�ĕ�^����̯m�e����Ԛ6��� �ڟ����bh��h� �i-�6v�\�n�|G�X\7��z��Kb�nc����Ĺg-����~�X	lXwb��D�8l���Ư��3N���Q ���3�0��cΠJlH�q{���;n�áU�0��[N#خ�O�f�z�i1���2�%k�ټ�ԟ�~��@�Q���^��a��:"����FzuY�dI�U"LX����"��Ȱ�'ͪV$�#ަ��y�����]cY�&��bk��ĺ��L�9��1����yݷyc5�K?�l�ƇH9�GpF�JiOoH\�n����e,W���>�!mZ��<*Lq[�Y��m�sF~w,��T�P���R�\��,=�0t��a���	b�����񠱐}��ӗD�*#�����_��Va3���vΉ�Д���L��M�R!�3��B���jM�R�*	jCZ_W����k�6��bR�qFaz���%úD���A\�x�"��Z�r$�b�,��&��"�����a��I�����T>����H�ޏ=CEA�;s���·gE^SY�ۥE�L7�wx�D��{	ؓ�.�Z� �?��нкC���*�5=��Ɗa|܏�\�E"��ȋ�� �_OT�Ԏ���%�l[&cj���!T5�)�"�bz��A;���3��wf�d�#�(a.G#ʩ2i�ڦS��
u9�#sf���.y*�nV�,hn�/�����.�
+gbVA~�veI9�9w���c-�+�5]���V���}���%W�o���!�cf�K5#�^#�ޓF�E��,�ذPE���~�>݈/]����'�!g�����H�Le�M��>RI�,7�2?��x�"�xC^z�B��Ø�[�͋t�_���%��i��:r�8��Q/�:ü�S˩��2�2�G�z��F�b���`˕�����Nzl&ea�����fm�i,��4��]��\��p,]O=;Xph�V���O��$�2C]�eǜ!d}E�ә2@�w7.�ޒWȣ�]pcc�laN߄�Jxm%>�Q=wպ���\�Q�}�QaALK�R�u��,4gQ���z����|`����k��7C8�k�������d��������V#}���E�$����J�dTX����um3�k��A=�#���&�v�{�K��»mIq6S��phI�"a�9@A,2���X��>X��6}����m"����G5N.��$ΚC�	��9�R��O���]yM7u�J��ه�wz�3-�$uW�0��N6@'�_�nVQ#a�˼���|����,�ޘ���<x������p��`HN	�D�g�Q�BHb�JN�KB� �{�؝R��S�/��e��SxB5�|F&<��,�>oU����Jk'5Ҡz8�Z�b�I�밒���.�L�L
�W�0}<"+���[������s����7�\�w�3\���Xz�-X����T��%m]�d�;Bh�2�޺��y<%���ߥw�	Qg7i'(.^5��o�Pف`��Y��{�)��ƾ�Rc�tb*�MO[�AP7�X���)�k�-�]]�+����k��ބ���l�%-�b��L}"�_:d��W�
 ��՘��瞫����C��<pS����r��F�>���,=��VAZ��YZ!` �Apt!�N���#�#�h4���k���F#�8����Ǉ���'j_wg��zK���gŦޟU�)��ࣆ��H������\�a�:>r��y��t��ށ���Ydy]�2�[�^_�NE��G��(�[j�F� �+VY�|��:�m�R?�	�Bǅ���b���W�N
�����O���%K��T���� ֶٚ�m�E�+EP�
�/L�#֎��4D�$�$�P�!RH���I&�МU����R[�}>��3rRƮ��d��5�ċ;������yq�Y{�ƅX��.Y������`d;� ��:N4�Ϭ�0Z�Iq*d�_�`�]�X�V���R=�|�y�'O2/�^�y���6�[��'W	�k��I�9���� b:J��J�c�L��4��06��,?�K<�!��eE9k���R���`}����XП[|��p��D_D}a�w��t��>5�I�z�c���rR�� �R�A�Ɇ�^��7�{�{� ֙mi�d:�i4�Ғ�fEau�Z�DT1/;v�%q�B�f���_�5�mk��޵��]i����?"�i��B����-�)������JAۭ~e�*#���7�G_���+��ik�G>v�0�\���L橐49ԙi�c�'����ݞ�r�����oƕC�;5?7X�� X���,�%��_Rn2�>�I��rx���!��<+,�I+�̶�%%%��^���/c3�\b�ަ����G	�"&"m��#�M��WN q={����;��D��<���5`N�YOi��T�8_�P��Ѱ>9e��8�qoP�{���G"�#��T��X˒��\�_��{�8p��ru+
�^�*���dV|�q���lxZ�	=��Æשo �����Zk���^ �3 ɀ�{�� g"��SB�=�NP��(�$Q��������)�ٟ1ݸ��l,oGFRu,���Ns�����ӫٽ3O�(�_aZ׀rҿSp��x�l��¾�t4�;|,C���]�m熃�hk�y�#cy�B�����!l��������|�%������n$���{@��A.��O�Mڠ-�;��۪������I>�M�cy
o��*}�����Y��:����]���l�Z�~1�e���4R��#�=���N�0	HN�C�Zh� 0�X�.��?�c���.2���NL̠�X`���7#�'����%����ʸ$�
C�<��bd`b @�U���r&�UF_�.����Q��	ώ��Fe˫�'矫r,a�����ܕ���t*�2�!�����eBY���J��$����Ǣ��;/��R��d��K"495�H��gP&m2�J��}�˹�1�z��M�I�=���{�H�G'hQ)�jO�`4r��.��U�Y�����h�Mn��ds78���r�����7WT���>kL jC�^Rb���1$�ʞz%M����ɯl� ʁ7���}#H�tv��tV��)䪕2��9�7{O�P;�L� ��/��T>1�R��)�"��_����Gn�Y�9��o�T��X=��"�OgQ�E�v� 	��|�QUr'�#L |��4Z��"�涁�3�)`@t-��G�Ե��Ҳ�P�fT-��jB�h�ˍk���/_���v��01Z���Yk,��ۍ���f�����X�%��C6ၢ�Y���QE�T����;�˃�!�����g��C��;�q?�_ȥ2����?J����	��́��.�"�r,Z#���Eں���=�+� �GL�>�(�ʲ� 	�??���(Sh��@v��4.���z�E��j���h	��S�K|�� ���V���W�B�� C�]w*=t?��p�O��˚(�Z�M�I�{��T�Q�	Iϑ����ca�����3L௢��k�?f�h���������k�ng'�R#ƙ�#��|^E�X�<��P�R4������R��*��cK����FѶB|}��4�a~ d�u����q%��8qz~	����V�슢���Qu�?��-V�ձIV�6�['�kMKN�A�~�T3�A�~漲�O�L3�G�򽪍JO(��֘�Z=<�]�\8����QN�q�)#U>��>���A}����l[��^l����Yl��?	�ƵFkfL [D��nd��}�$pV�.3���N;����&$�^��~/���7��7�
��Zk�۩5n*�l��{��͖q%�Z�Q~�!��L�W�c�w��&Bs��8/ys�b�vn�F�DVζ��*:p��ɖ�@K�2xc{�|��f�8��?�'9��/�N��6֪o-�7?�D�%2������]C�K]ݟy��9_n�)͞nU��䊇.�9Ua����q4�zG���:=�5�~i߲~_FXG�@;[pD2e��3�7^IJS�v�I�?r���x�zncC
�������VK0�|�dKw��-H�����p���'�j�"�W8����	O('�y�rr���<������=wҘQ�,�M,R}.��g+i� U�x���#j��FC�"Й�z�Qf�k�Zf�.�ٷb\5��DQ�����C̃�V��4��E2�[�w��:됟��H�I��U���{#�����:?��p�<���̂�����)#�:��	��������o�P�9��/N�����v��a��n6�	��v�ӈ��O�Ӓ�c5���Sн��=�[�4�4�J9�g�1����C�$��o�6{�%h�8��Ͷ:G���M��x&��Ȝ�<hO���n`� OC
3���!�L��*��8���\�g�CM7��W����,̢A.�0��켶��Z?��b�'��ɩT�s\�Μ��_b$�����	�=������>��a�r�&ںY뗆mߗ
?JQ�U,���G��Bn`8G���#��*�C[��gn���4�؉�I'�>�"��v��/�g*�^e�Cn8�������<b?�	�dg��w���F�@��\Y�޳7�	M/�-�xú05F
ϧ1;�lݘgk\D���_ �"{�1T#H6�]����&n����y��׷��(�3��y�v}!����K!C����/�in�Ih � |5������`#�NNE�������ڝ�FɇJ�s�V�P�Hk�$�B��0>�ݧm�5�ߵ��V
�d8~[79�(B��C�� �쐟G��u���	b7�}�vbA�Ku�T�@ǳi�H�e�����c&���g�s��95�'�u�C�9&��X�K5� %�Ղ��\7] �d%F��3�����[���1�ZS�|��Q�����~2~�����"�x�=ʟ�rI�B��=8s󉊼
<�5�M�i���68�����q��8��$�;X!T�y�v������Y��6���y��]7�郁�qF�;h1�g]P�y[=�j��4̡�ΊPw��	�|A �F�>/��=��E�� 6s�:�'�q�58����t���y@�l��&�z[���4�C{���4t��voW�i�s�u#ALz�$}ɬ.�!���kFK��쵮dʋ2c��[!�~݄�EkW�bI�g���k���٦��N&d́��W�Y�m�\��۞JO!<��%�c R�3x=B2��Q/�j+��'ǚ��f#���߈lh����R�A`����
-Aql�_<�����ģ��;Ґ�F�i��+�&؃CR�FlV��� i�&|� �'1��1�&F8�><}m� 	#�齐��um�,\�ʜ=����k���ѱ6�\�Pq��ptG�,� �n�g����]�JFt�M��KkT�5=������P�����v��z]�R~�9����o<��fG.���j.�dZ�rǗ�ҧ��\�<2x�>r�ϗ�{��9ί�#$M�N�:牛���#��Y=bѐ]���&4yO��I���S |'WN�t=�X�������v���M�������^���o^d�j��&���y��b%	��^����VEN�oFI��7�t�K3sI��m������K�J�c�B;��}�$?��;��=��h�ſG���&\T�䮱l0d?�9D�,#hUQ�9yI�(ڋ(�C��U�pܥX볙�� �P�� �A��_�CBA�+m*���T\�(Q��e%_HД zT���Q��7��_�`]03.RY����2=���(x݋���깟��韙�\�ׇ�|�=��C�J��F8a�6I��bC ��4Z���&Y�{��L���`s.��S�0�S�0���[Bu��/P: :C�s��~�i�MB�n�{��
8n��B�K��̧��2���6��Q�q4)�8*��+��yY���te\#�f����1�n�m�e� �<��P�M��xb�v�S�i�@����Yt(�܃���"�#����F,TY���x�4����~���ŉ�=��m��f��<��M90ܶ�}!aR,ݗ>W������Y0�/4�ŨES!���bĽ3�Jw΄�<z#O��׬�Q$N��ƹO��!�}6?9��o�hq�����m�`�!~rm8)�:K
T� nԸ.)J�9�4N�Ş�f�1:O��:GfS�V��U���YCڛ_v-6r�cՉ��H�C����r�� t�f�^
���S�탧��ݚbn�{�bӟ������;(J����>��
�}��w��j�w���`��~��r_-a$Y���Qr����QտWM�Rh�����OM=�Q�'E��d��!h����aݚ.�����#��{RhIՒ 9��PHD�
娰�M<dH���&�����rT>�zͳ��/q~�y�?X�g8W@�3��mV�{��I�|����9�x�̿%=���voNq���ɧ[熟p ��ṿI5��tn]���9��G|@7��@�h���$����d_�s:�
�S���
�S�/"��E��:v<|0�j7;o!鬻���;����CgB"�ŚVTg��h <��=��?�9�N`=_��?��=׎P��4���cAe��2,V��M��pr��u�lE^�@���n<&���I��)g�As�"p��no���+q�d����u�w0f�D���[lXA`���(|���h����ٝ-,�e�Hݎ�v�s���1����S�C���(��Ė�ɝ﹤D[1ͮ1�D&��A���K���O4���F��VBoEf��}��Z��L���	R�&d�B��=P	t��Y�u��ȥ������c��t@��YС�)�mì�x)|���+��nƝb��%R:�$5� �'�d�������c����tN��wG��6nS�f�f��z�*��K{��&J"(�4�$�C��׶"�6o�?�|�|�o�Gx�5�7�cֶ��
���1k�a�M3�ýBO�s}���8�HKaF�.�Q쿒��M0�����h��E�שy�����N��7�4z%}qY��.�^�#�_��"Y�KEgz
3US�&�9v�,��ª� ?�!���
��:�?8!� y��l-���5��fs��I����Dm�B��Y1�@k#TI�+��C���L*	3˰J�G8�j�ۀю��A�Py�Hg���vv���>���~�늉�.;D �E0�>l3 �>��l��+����A�:Yݢ��E�S#)	4��@��q��vPf��6�K�wSi�Q�E�$�p��߾���O�5��zW޽1`�%Kt�g�Ӹe���n�孱"��A��ybk��p ˽_I��e���?-�͏ ��=��׍�h�.�����;?Y�p|�8�CG��$�}�{��N-������N��Q�L��!H��լ��ϧK�
��ӀH�w���
u1mi�b]/�f��#i��5( �
1�X�`��k2-����/�0xV���%E�gc��}��=06m��ޫ�~�|�ȁ{v�� ;Fԧ�*8��_���q;~�l�qѴ>4^/I��B��Xt��	lO��wӒ.�#�;�6��ܴ�g��}��}�b������l��l�G����^���u�$�]����5J:�w�o���o����E\�����@�:��g�W�eUC��5���8�h:������12=��CDl�J�N��3<3��I�e��RV2�Z�Pc�v��w�	���3��`�b�pʼ!�`.ooN�5p7�钩ɯd����2�kN]ǵ�C:�3p��L��i����I
����VIa�]]��K��.~10Ҽ���a0KS2:-��[� �Y"��	lϻi���$��sZ7z��ǿZ0$.4ɨ��@�#]S7�7N�i��݊�O,/��d���Ϙ�G7@k8k��4Hl�p�ٱaR/b�F��nw04Ln>�����d�;�2[���:q� ��7)FC��2�j��327:����B"t�X���u�8E�Ⲩ]�n0Y���V�Bǥ9�����W�H��0�"Ķ-�I��7ȼ-�䋢A7:Ǉ�(�x�;�o��K,ȉ�aEX��	�����"�Fd�%��ML��K����z����a�H0/���M�r�9�8Q�跞kn!F#r��熈�׿�����1�Q8�J7��}r��-�F���9#������Av&[���l|��o=p^�J����C!J��k
��N�G���	ls�&��թ�;������˞�ۇ�z<��ڿ�����F���"~��C{>�`����	����}���' s�	\� ��GjLO��y�)�إb�Ϫ.ޞժ�O���NϕZ5i	���m��ɭKzVt�O�.�9�Y��J��5R�ʉ�KX'���-%�z�;C.zQ����t�H^�����s���6]i�Y�o���X�%��s 3>5,��]�4�7.uT��e&��TPblG	���ࢠ
�+4���nD��ǚK�V(�,1l7���3�I`{��¯�`���0�T�v��M��;Em��H�~�j����ac�������P�ݶ{���Zt��2�鷟S��Yʡ�y���Z��%�	+����I�Zٸ���
	WΚR�w3I�>#����='�t�gacvb�j��g+�(h5���I��Q�Q���v��3���������Z���F	�?gQQq齲?�%B�Fg�:qz,�����Y��E�����c���-mݥ�ª��>:S�c<������Knʧ�1�h,mm��K䦟���Q�S�KIσ��V$�my������	�z����m/�����U�Y<�S��ll�dl���a����;�H�U���n�5�"}Sb��-����R�2.�G���רc�����\Y���ܖ�}�׍�����K4bB5X�u� m�����o��c?w_���l�� z��=��������%��D� ��q�\�f�c&�s ��E�߯n��D	��SA���w%iā���{K�&�??X\�>�����}v��g�������U�s�LM:x4j�U{���H�q�EG$�K�:k#5~j���e�Ĵ�!�uzJN�48%N,��(H�E4(�<R7zT�DV?�8�h�n8	��@5��z"@���_���{ôy4�=��B,�]0��=��uLߧj�Xzw+�@�)f�g�aC�BO �&wXUv���I9�cP] eX��(�][ɤY���Ud�@�'��*�\�.�v�%J�}�$7PJd��9��A�ށ�A�D<)���?�JgA�N{E5l*t�d�]��=�������]���%�%�j#�c}����	��'{�Z��Sށ)�af}A����c�z@}~��P��,�wFn��/]-!�o�dy���?��Z��ϜT]�x����~1ݍ&3�I�h�@��)ɐ!Ë�XZ!!���<}b���(x�~���$8��ak�C}�m`�$E͑>�M�2ڎ�Ϧت��D��N�BI�V���&�f�$�?�M�]��8��:���k1y�rq�PTq�[�y� _����^������3�#$�S_�w#�&���aP6�씇j��Y�G�U�0����L���H���q���+�{�v��
]��;!h�NRψ�D	�֧F9�?9�9K)�!���q��*i����=�x�#����7���86ڱ�U�0j�E��m籨��W-G���(���;!q��m��T�7l���ٸ�*��	��&�~hº5t\SZ�?�]Q�LO�O��n��/�/���d��N�ؘ����Z�0��L�	�A�3w��Q���
��_ij�q�}=��@i~}�����t-��u�k�DSv�&Q��D�BA �ך����z>�y%�f�iM�}B�/���
]��.p2��tR���Ը��l�E�Oy�����Ay8��ϯ%���n��h�쓦k�B��@���B"ZL
5�b�kC$+���
)��������7?i�NWE/>nω�	j+(lClR?�E��:f�{ F�x�g����rW^�%v0�"������]y�� `�,�]�%���-��A0<DՎUبaX"���(�i_�) ��� 2U{��qYj�%�՗B����0�S�e�-��7�jq��[�SY��݀9�ي���)�a�3=���S�;�SƲ)\�%̷b�'+��=E�I~T��,��*6�O�h�]�OoB��0�a����+������=Lkp�$����T-�����k:�q�'(�H��+�g"*���XӢ5Ě;Gs�.����l�or��R��o�\nD�\Z�mm`��j����D���& !P�����8$�X��CO:��=�;��<#~�L4C&��Cg�L!3̥2��D�/�S����R~�f�V��֥��돝�ûA��%7�?������B�3Y�*o�d���%��k��"p��hIr%����HL��W�ٷG�p�\|���m�����H����v�=p8�����%�U?��������#�eiW+9]�8\�}Q;�1O�� Yu����y=�`�}�>l��ŏ�z�S��q&j�&�F��b������X�u84,��:lξ�
�B�Y���e'NF�ѣ3N�"��4��"�a�ū����v��p/��)}��'
�����C�� ���5������ː��&�>wT �ݑ�b��NM���ӦS����ʛ�����ch��p�D ��V
�j2`�x:�T��3��5��<x��Q�����#��~C%�P ��W�"I���C�tD�����������Y�2��#���wM���!^���;�'�J}��ir��6�O�)05�����v=%ejy����1��;ڷ�r����Cˀ%�R���O�{S�@2p�3G��:H�~y+P���XE�c�ץ3��vGq�y��:�h��F�����M�,	.��F_[�M��67����Z~6��d �Nu|�"��O~�\�d���]T�<dL,�t���L[�J�#���~�������[N�ͼ�6O!����W�Bn�\Wj�M^���c>/��̘=y`����3�J���X�9~0\�`bkD>����a��g��ӯ�̂�v�w��X�B��P��"*�&������mbn	��&�w�f|@���㇑f�a���i��g���m@��}~R�]�0/�kL�@������.����!�rC�*��U.�����K ��;�F���
��䶍���_�r��O�Om�-���\����u!el�$-Y��`,AbG��v����k�+*�7܃���n~Q�rk���j��>*�%���J���#h1l��DNt��Q�����P@O�����o���ǉ�Ý7�(�J�r�!�\��6� ��P���V�;B�����+��-6d 5Pߊ�f��bRr��p����>-7�[���^�ӥ���:ƶ`�|��Uź(��"L��İ�1x�fR�1��è�X�HHI��9E���F�2��qvwjfq��!�Z���".�I�DB%���J���nJ�`"j�Q�z����Y	��{+�^g5���d�eǉ�*S�Àu>�e�J��Sd����s�đ%ڨn�os�
0��E���a��c��pq9De�j0�53��έ�	r�nRA�0��W�YO������aCh�@#��A�W�yp��[L��S-����f�ă���:Ë�s%�T쇲�& �?/�~�+gwz��W�`��M������(pE���b��S+�O3@p蹘 jT};P)��g*�*w��{Y���5E��[hӔZ$�d�X���,p�S�s�I�/���z3Ka��{m��S���s���x�&Oj���T!(�~�m2wa��%8}Aa�1]�F�B�#��d��n�=�$��Di���w��-r/�ećsE�$0?vvv���Ж���i�vZ �Q��C��_Y��'V�����p���T*���]����
�Rs1@���L��>�h��x�< o��-�.o�;8�Eyɀl�i��I�i�@'(<�ν=Vs#�/LБ�n	^�A���۶ oJ �WM͹���&�âd3�8nV�קUk���Q��2�k�K>��{���ף }�#���CU���K&��
��~&ڊ1��A��~�]���JO7@�zrG6��a�H�roN�`�ml���m���Hx���5���}�=�K�<�;H��x���P�����n�F�x����E9D*	nv�߸�7�_��g�P5[�X��6�2\��3�g�ې��o>��{�)M��[|3_�뢣c~�)C������ p�Go����C3�Iڭs݅4�G��Zѽ���m��զ���� �I+���pJ̓2����Y9K��$����vXZ�gCbh3Jx�`M��|z�o��<�~��-x���f�dz-���5�ƍ�*�Q�f_\�G�L^�ί����g��a.�B��9�����N�yٌ�(2�9�ٵ�
�$��݆sJ�X��g�ah�����wk�'8��'O���~�(.�%�W�:� �u�싷�e+�<=�a�������z'OH�&��<F�?��L���F�q�|�Wo���2�Ͽ�:��t���|"�2 56���y�_�U� ������Xi+��Ӽ�J��w�u>^{Q���uU=r�ETRW��Zl2��J\.������VU��_Ol���-�H�-j�í���@�0��<�魹��;QS�f���1|�5���hÎݿ��9��A���`@��u;1WHd�y������ԈF5~<L�u����i�'�D���}�e�,`��o��9RL-5V�ΰ�:&o�������nzT�i��s^�L�&��GL�NX�9���V��1gH3p�l:��X�a�:^/�oژ�nFD��b�^�\c�M�z9��F��������n�D"��C���l�n��7o�!p�PI���;��?��mL*^f�3MtC�E5�K�KH+���̐ ��E�z��-�TI3�ʥ�M�_�d�~*���oL�Oc�ĉ���l&�N�<ș���
2@̒��dK�C|�2��*�X{��V5q�aj��fw8�!I0&�u9>졺�Sn)�*���J�����튴v�`��JH��~+�Ý#�F���:��nE�=m
�ҵM�ږ�0���T�]?��h+)��fl����l��m��ý��,���<N�c�=�s�Z������O+g�;�W��-'P���1h��_~�'�Ó������� �9M ±��!d�[�͇~��e��?�D�}_� �t!l6�[l�7�F���(�N��;�I�j��仃����$��ĝ�_�� y1��S�z@ �PE��!q�K�i��tPnN�H#O3KL�̉6IG����eH����GҐ)��ֻ���'4�1TR}�R�Տ�x����q�-��ï,�CQ{E��*�7$-,0��;;4zQJd[!Dg���m b�j�dҊ
U5d0��+�u�qy�ܲTw�NF=�0��۵�S��j���6\�JNM!)1Sw���-�����L�?�蕑��8�-�u��\��S}{�O���+��\�����\�0w&7y%4�u��|�&��.�	"b��)���	�l_�w��*�qW�ƻ.�b+�-8��M�lkT0�lS:�,�fj����Q�, �ä
��AHz����Z�iF��h	��cq�\�qC���u�NrkWk[IR�͵�P���#�fF�$�z`l/�D�-ON�Wy���07 �BA����s�!�ss,���4X�.[�;����bE�n����O^0#�d�3��$�?�3d?6Y��a �Acb�'��j��];i3_Ǳ@��F����o!<�,����m��տ.�k�>ḻ����w`d����[i���q�Tł�P
e���KH�ƒf$�'.��j�"�ҳZ[Z	�̈	+�^?A�.L�u�)_�ɼk��n�Ƴ� Q�S?���G��=�񧟞�{��}�.f	\��[/��L�j	Q�G���ǝ�QK�,^u��l2<?�6#ƜNЍ �㢟�-�����iZ7o=�`�D_�ڥ,� εb�;M�]uN��?�Sޱ0NmXp2���g�U`�{UK(m�sBu�?T��ʭ���И��qşVXh�P�n�bm�G&E~X�fx�w��k�qtd�ĪE6��΅��˂Ό(&G��C$�������:��A�`�ߝ�AHv��73�?�ѾωĭK�q�ԘPq�j�k 7>����C��(ru�˪�u9G{HV����B�;�EC�f.=2�4HkDN���*�'����eD����#7�U�I���$����쉰Y���f�����M�y/eA	Q�o������3�Q;j�<AJ{��|�YV�Ę~�ѫ������J4�E��eN-8@\&��jU>�	=�+�E�)���u
/�٪��ҭ�
v��y�s��� '�T�ҝUV(��L�w�R�I���aJa�t�*�_�͉��V�R��E��Xl`�Z�:>�ދ-
jc,�C�&��-��#����v��D���%2Z��h#Q�E	�qmO�&�˦:�\�Fߍ��#��\�~Q�D�:L�]d���,�>�P�����H��1۽S�f�=fX�e/��Ddz�����\���|e>��E}9�f�<fGU�<��G^R|D�:H)w��u]\���J]͛o�t��.1�H�����9h�~���U�!͟�?j4n����'�xH]���%�wb�.L�bN9�8�$���q��Q�E��N2 ����[[��3^A޼fu(U�kujm�B�{�l?>��o��9����HW&/2��G�;\�`�Д+{�F$j���.�JP2���p6M�	�4<���<���<����Z��{�=�e.�b�"�+Ӣ
b0en�7uF�������*���R��)8�Dsi����I�6'����W�7:���@�G�K"B\�*|+tIo��9B܎��Ә���N2!�c�F��p����1ٳ$@�!�Tl�1U�2�G�>�$l0ߐ_+h�Q&��/F
�>2����+�hsz����!�
�-��vB9K_n�a�J��3=���%u����~T]����>��%��HW6|�u[���i�P��p�VUJ\��0�.x��4yr�v�b^-�V-��f~ӂr[�î 5F��>o }��K�.��>59���X�/������;0��&�3e,��Y}Sq����h��V����<9:d�=�f�W'������L���3���H� �w��l
��glq�x�Lyو��"��g�W�*�����xG�����Y@��nΰ 0	O�� ��	�^0�y�7����l����-s�����5�S��r�0��0���[�6�.��J��XYL����s"�����{<��WBSh�:a�P�b����Q+X��?��i6����t�4�N�.D���7��:��~4�ЁM2�3c7į7�8��;����u��yjq����C��ӎ���˵Z��'�7�S""���WU9~�P�H�PU`gH-C+�����qtu˼���SX�+���� s���x�2�H�c�,�?��k�Κ�ym�hJ���손�jَ2�#���1D�ku��/.w�]�ru��Ms�*������_A�Y�E��M�Wߟ��s�~6<�v��'���#|:v^F�Z?������^%�(!(L�[�8yo@N��P��i"��>~��K��Z����X��8{� ���Q\���{U螕T5c>�&!� ���Yc�9�N�=Nk�l�/�������x��k��������%��٥�鿁dP����AK�����v�k\�8�F%6bn0f��{���1h��'ox�6��1��Z+�n��㨛��|�����/��?�s1��H쵩���(��g���pSڄ=(�vn�$0^˪�\�V�-��W~I���vtX�2��k;^Q,��iS������<qQ�Ȍ�~��S��D'����!��rD��b��
Z�z���b�	��m���%>��Q�O� ��u;�ǁ%؎�H����_Ҿ��Y8H��8��$�dV���F_y'�q�J����ݸ'a���4>��h��X�7��n��Cߚ��=Q��� (�R*{%��?��bc��YR�����(�F�y����a�V�<T~�}�.{�J��ګ�2�(ѝ�@�,"ٗH622����;�p��- 5�h�9��L>A1HG;,H�t�s����4"��K�p�T0�VjW�@3�L���L�χД� ����?�V	%7ՌR��9'��V��_��}���]pߥc n�uhWYt�Ytzl:�@f����F���ɯ��|���YԵ��A����-r�����c��{�β�|�F�h��$p��{)��?���+G,��h�ŭ24`��OV��jUA:���ɪ������!�W�O����u�&`��H|O�"ف6�S<���^���ƽ!��Oc���uT<)��;���x᳆���y�:�Hd��M�8V9��mC 
��-��Мp��?�`%�4�n¥R8U6d�8�;�EH�Gg���]�(E� y0�>�C� �S�h,\�{�̓�$^̐O̔G,�Bj�+P��_+��B[	��Г�~��Ҿ&F��`�)'����ў}p�e���/=S�u�~$I�.aƏ��)���\o<�KtL�ɀǧ�ofm�����g\��%�3��u��O�b�M��Eo����������|̞�3�<p�>���ۯ3���b��,ɴ����L�87�ݎ�1+� ���f�{,z�梂\�NAU��=��ن��8q׆��W�Φ�C-���>�LtXM��Ws�Wի׎����9T�>V0�۲$巏tt�?���T�Xq�:v�}1�~� (�	���I��Z\�o��������/荰jG(|�16\!Ӏ�<�UKdH��%:[����f`� !�D�jzo�?>����~�j��6&�uDe:R�$�{���=����9+��19U"��Vτ����w.�/
�i�$.8���1`7K��4�o�\'���au�����]�䌎�*5D�A�����Z��N�g�o�bJ�.��1��l�;f_��1�ep��>nz�ƻ��N(��v��Gp٧ᛔl#Lzq��7s�=U��rkCu�Y8s�㏑����X�-�>u{[��[d�G��~�몡�ęa�����^�y���x�M 3E\V���8��
T������3ɯ�_�UX�+����q��qj�C+g�( ��J̙Ol���pQ��xF�s�A��|��E�H̽_m�<�jw��tx��� 7�^�|�T��P��Qz�{�@~@r�pc����[d�HΧgۄ��=ʜ�&�������L.���7�N��S0
��G��7j	A�9��fv��¦w��"w�J/_��u���!C��R������D�c�/����-����:��Xz}�4�0J��d����K�����4��s� ����_����d��dr�j��8,��ef]�:K��iҴ�S�{�p��a�?����K��Nm�8�q�H�V)��4�1L3T��a猎�Bwe�6�ނ7Є����)v��E"ܳ�y� �w��m5��9�Q>Z�6s�F��ɚfW\�>���`�O�X���V��(>c�Ϟ�	mȴ4�1"o�o����N	��k�5 !�I �ދ!�y��
P�=��)F��R�ʹK�]?k�_�����7�n��w���+�*��ha�ab͆r��i��g�l��o/AV����/eڽkb�i������]Ո���x�d�}"�X���9����sK=�Ĉ�%p�*���>������U���u��k��)�m��aQ{�6��s�؁4��N�����m�;����/ �F�zC�NH��D`:�)�?�o�N��̉ ˔��8���[�v�[��B����2�,��ogȚ�a��]\���a+#G�v6�"���
p#�Z���|#A�%�D�T�|��z|���O�p6m��Zj�#j��q�8�wV��j5�����m6��\8'��4�K�|7b6�(��|���vL�6�A��)�( t�Y��gM�voX9ʓ����N�Z��F������/3�"wZ�
�����?�ύ�jឌ� k<`\�N`�W5.�cTh�~��5��t�V>N`rgU����3�/6g'��_(0Sf�J���;��j?*�R�yU��^��02��f��pH��o%��g��X��A0蝋�u�j�A�#f�����-]�h���ȋ]�|�
�:ƪc��(�&���2�$���{~�u��hK��v��_�&�����X(�|W�#Y��I蹯okv��С�V�aNMA�]�r��~tȐB��:�gC��
��P~Q�6�ԫ�>�y��)�z)�=o��a0��*V�ps�fI��_����K�I�U:G@:��~������y��R�QJ�u2G���O9~+ܒ��4�n�+�lC2��]�5d���l�0�o�N�U,��T��\qK��o"Nqy���z��f��	�����؊�Ko��by0e�"6P��ߨ=7E�f�_iD���|#,��J���ͩ�+)�!N%��f\!}ZAV_ �"�x��}b�0��0@;P���é�N׀g��o���|�Z1E����VΉ$�t���ˎ�r�jD&��bzj!�8�)�K�[+��#1��h�+ Sn��Z�3��@Bu�u&����w�w��B�,ٮ)�+�ǊQ|<�-<�-F����/�S��V'Z���<(�5<%՝$�6H���D��/�j���������z��/��`�c&1�Y܄�L*�K��h&�)7�5y� KB7�WEE�`|�k��(����Kq[��j�wCopZ�i�X�>ՇrZ=QV���BS򺼁<B<6��U���̖�{wRN��p���3[Y�4L%��{����U86�Kn\c��fѣ��)��;ѳ�u� �҆Q��,�Q9��E���w���v��ӊ��m�d����[��NZpg�1��'N�-�U�=k�3���:'

�� ��3L��HI��J��C�ֈ�2ٮ�{+��*�:�C`�ch�H����������S@/��De�W��H��VG���Q<��@|�i{g�,�;<�vg���*��@���;��(��d9<�cF�gr�;��&�Ef��(�8� 6W��:A;v��
�խԏb��˞�
y���&H�-�b�xeƔC?rR9{\��iϷ�[r��.{Q�)��gvb�!9����sN���4y�f�X�C�b9f���Q@b���Z�A(�]�ãI��ے,)U����\�r���ǆ�)�@�b?S�)��9|X�5g����1&~�඘wzS�8A�(���E|ȇ8�q��0��c�&���.f0�3c����PUH�l�_�1kr��d8S�w,�@���J.��q��A�W�,d�4�ƻIi�:�aP{d���cY՞������oש[X����G�ϊ�_x�Y�� K�'�\��S��\�v��>�62��V�Q͏�y8aMzï�m��(k]Ǭ紐�Z����f:h3�W��ә�D0�f+nGE���p*�������{�Kz���'픴�y�D�fOQ��׊�
��7��i�y���x��G�~B�^�_M^[���3����	8�$C��%�.��5K�x�٘���Ąj����U��~�6'�7����Ѳ�|���A��X��i9d�頋̠�ڄGő��{!�[�\v���QU�{�9@d=��E�TG�W��0�T��+�?��f���F� �4�w���bz�ĺubX��:}�I���
�/֗u��鲨q&fG�'\#3�7��jO�C������;���\�N��"�$� ���i�U���Nʋ�I��%Q�N�"Q�77��Xh�X�F^y���M�i��'�Ղ^�.�M���P~ 
a�uMٰ%>=���=	�u_Q����6�����𜵈�N���9�������{���]����6~ʞ��gk������(��(&�7T�O�q���ƫ�c��v�FX&)�^�nK��/sS�ת��k�S�H�	G�
�	��9[^͍)E{M���)\�ά!'����Vt�(g��!�N��9��ϼ,#�3�O�[G�\�b��]5b���#<QK�i�@���0q�f��ľ�M'�O"D�*+�j�)(�k6r �6�1� ��$�X��slV/x��9�x���Иխ��a�@	 �}�y쑡" ��R�R�]����;�h2�fb&`�Ū���� }����v��ѧ!/0$��p�a�|�]���#i�Ӡ��U?D�+=�	��oj�|�'�r���R��-� �\$�5_��,�P��vN8��%��i�^lrժ�Ҍod�*)'+�?K᧴Gn�e�VoQ��Ħ	�ud��Oq��M(�-;��%,�&�`�k�p_Ig��=���ǎb�3���� H<52FB�3��WH��*��̢�z1�,se���L���/�����K~�$^������)#��SZ��	�[��[E@U�d�.a�~���]�i�,�[���Vo�'��w$�^��N[��a�p��Uy�yM��0PN0�Cv��'��;"2Z�Wq7�Ѧ��tE�Qф%�V�?�"��[���{����{�v
E�s@94�VϒK ��O�Ay�l9?t��~���6LJ@��C���aA����e�_�˄d$o�T�v� F�1��ӿ��ڳ���ٝ!^YU�U(�����f��H}�f�	�hUβH)ǒ���z[ݛ��"���=u[T��P�"�(�tyh_.%��NS'��`X4�o��Hz�����+��5�q���8��^,������|�6 +s���iD�\c���Q2 �3��6L���FV�dR�}���&k	-Lޠ��ũ�H�V�6��V��c�ԵLj~ٗ��'E��ԚI��zd��k8]�%AZ��~z�si�B�b��l
;�\�F`.h2��5g�e{�=�I�	�����w�+Q��lP�$2�>�0fh!�^u?���p?Ȝ�t���+:���|� +��{m�8�?x(�(Ve zLR�'ev,�_�j�rυ慉%ҹ�����ݥ�(~�픀h�L���|��yNF����4�+-X�G�C���d��c�ϐj�r�*��۾g,Uo~�G�qTd�x��͹���*ǡTK���kx+�h�`9�p�Н����S����S_��R��(鏵e�	��N��OCR-�LU?稙��P�����_{n���M�r^0��1\��}ޮD>t�A�|��K�X�S��Bf#����eP1�+a�طP5�� P$Z��R�x`��k����6��P!K@��j0�h�������m0]��xο#E6J��A/C{���B���;O�ނ�Uz�ޜ�l���~�t��U�p�BR���-ݳu�����尓8Y̗kۓD[�j��.&��ව����k��4������xT �u-���[I��
mhq^����> #��>>��a2t�bH*ܰ@��;��W<����|R��Ӡ_!��1�"a~�7cd��×�Ĭ5�y��r�F4k:C�5�Tғ8p]zJ(��9Ka���h�ַ�!G�N�b_ۭ���v�R��¤d�hl�H�����A��?6��4^���k����0��~]�
��/&��ജ|�ϝ؞���_�P����-�	�'SAaE\M�̖X:LH�Up+��x4�� 7'�'`s�@�k��]�+�L(Y���$ybo*1J��ZZW�$q;Lv�?͖hO�
d�����r���O�Lٖz�+���w��e����~�yY䱨�MO+�=o6�4�Q;�o������"��s?���=i�R/f	�Z��K�N=��=��N��Z`Ma\��yl�]��F�0�V�N��Ջ��f4F�fV�9���NN��D�/D�?e�# �e���Č?&IE���bӳ1AO���t]��+QDr�m��b���sQ�!���K�z��̱K�v~�xrspH�5��`� ���s �E+�4���%�O
� OOdr���� �щPt�a6[�91���b1%���` �Z����
J@�j����*o�/���}��Q��٩����ZgHLT�$u(y�V�a�>9���^�FH�",��r
�Y�6���҈������*x�U�Gl���N��I���/�+��>Q#C��nEh��ց:��?���:sq�;�����tp�,�@�(w��|�_��ޚl<4��к��~RH���U�b-�pl�͊<ٖ;>.��.�QL+�?�};��kqs�<JA�c��ӈ�9���,��Ԍ�ͺ�W�@ݘ�k2�� s�����9�A%�S�V;�i�\#�,�����3�5���Q�D��$�M���;֩/�r��
�E�4�G���~Z�4ݧ�s�[��dh�ȭ��0x��:�2T����b�K�h��š:��=��;�����|Od��n�R��j}?�5��|�j�l]u�l}i�~�1L ��4����W0Rk|��
��9�;#�*��+��{�M]�[�
��f=&�ȅqڤP�?�fa�mFp�M�ֻ�i�9���'�q�*��p�إ�0"�c�f$J����j�E��9@��ү���;��7ς�0M(-�5�"�+����>�8��_6Ct�w�e~�sR���[�u�[k%t��!�p� �7�j��a�����#]+�u���J@���s��	�Η.ۃ�k��Y���_�`I�9���ځH�yPC�jl=�rX%/�x���C�\ Jo<]�Y��ˠ*���pnY�G0�+ ��A�z���\=�8.�c�Ș�B�֮۝���B��5������J�K�
ľ,`WX���OF�����T��f��qC������Q�:���!Q1��FD��,%��%Dپs�~?*��ށGc=e�M:asۥ�]���w��Wͻ)~����̗"
M�-9�߰m(d��p���g�Y�MK2xx{v�Lָ�?�=�T�E�-�\fޘa�!Q�� :c�oC]�C<Jz��mJ��]��M82��c�W���ѱ�@-����E�ٓF�W��G��xrj(�@,¤ҐdM�h�s��=��nx\U��6�����	�PZv�d��Ž�?�K�Y)rb�ڟ�-y����3�)n���Ȋ��Lo4�;
��6)�(����W��!;!=���(�\\켈��IB����!�[�̊��؁�Ͳ<}��^@(}T��~�/�p �����&� J���e���L!7�Od�r��>����S�T�HŊ&q�S^���W?�?��1U��_@*�=��(),#��!�Sn�ᦝi0} �S�!dru+��$:mǆ�U��8���J��kOO�C J��N��
�H�����d��Ȑm��7Ç�~�Zi4b~�s�:)F�g���#�$=��|N�����ry�9Y�f$�;J�:��j���n���^��"s3���w�������3�$���a�?d7��'�`qz�5�pʥ�ʤxD�B��k�4�+o��X彬Pz~�,�s��k�o����Q\�k�š�PhW�-���C���Ai�NK>�2�5�brEYp�!7Zh�Y�ȉ!JP0����#�������r�P��m�Κ'96H���}���w�R���K���F!F�ފl�B؃�x��(0�yƚB�
�>c��4�ݼ�_/ǔb��d��j���$N��x��R*SBU}%@ϧ[^ l��3���N<�橏��ފom�/�lA��p���ױ�<��?0\/g�<ύ��Qrq^88�/�1����ELUټ4�y�A�V95F+4Îb�mŃp�p���������ߢ�>x\�[]�W��!f�E/�r�yч(��	�E��MPcO��-��D`26��b�u��G����q����L��#o(œtI^t�w�I+��V�z�
h؉8*�
���~�r;�G���O$�I�		5hnY�S���]뜛���V�q��ѹE�![��*Z�\)ӂ^���A�S�M9���4��d<�K�E�}�h�)�kuy!9�8��in�{Pޗ��L�P5�x��� ��u�J���Ӽ*�����cE~��Kr��9���e$�Ⱥ�$I&a!��ch�tY�0u���P�{"����NK�P:�)]�~�ػ`�wu<�`y%��q�_�^ۀ ��t�I�b[���!�)e,���#"�/~�k�-�����&��HG��$�����9oGp�������/��}�#���	�z�5���fj�f��H��$�9�At��~!>IV-|��+�V��?ⱈ	`��(��e��uK�+�V>�(��z=+{������1$���l�q4���ǇN�d#?g�~�v�3�Ҡ%by��2	����;ί/�)6�ĵ�	����V�m:��,a��.�e�%kҵ�[���	I-����г������_ J��G��䬽*�(}�?TKRB��`C�f�;�6O܅t��G���?7tx�h.?���fD�6܊���w1�b��4�w�𳎆Y�� �������_b E��J�Q!q�_	����H�M��ƸQ%3s�?�+?�U��U
�`���h�Z"��Q�lԩC*�[_L*���x�%,x@�źN�`�p�����pGrޛ@�Jiw�D1�Z-�U
}x�Vi_��W�v�_o�F'�]����t�c�NC�m��u���Nu"�N:uv�PF�K����$�^pF�SO�	�^v�+GGpj-��Z�a8�Ҽ������I=^ӈ��f���`�.�a;Z��Ǝx��(%�Y���������Cϝ��~��s��`�U�8D�p
^#V`�O��w�h"df.Nb������wȻO=�R>�n�q�}�k˪w�O��1��v��Wc���%�ul����bQC,���:��CZ��Tb��U��E����w�!��
H��<.�Q``�ޡTFyF�9�.H;�9�~�C�v�x,ݱ�g����tV�r���?*�&����b`��ף)�Y��9�7B��]Ap�h�C��� ��ϝ�Q�D��3���{zz��9[����=3<�BP*��`|��u0ԁ;<��r��b�q
��t|v���ő���I�b=��W���������@��(��bXO���L.D�����&��/����z�0i���M�F�l��$���!�[I���M8�:�!
���ȇ���,���動�����*�]��c��^�:��x�[= �Ȕ���a$D��s5�4�Y��g��_Fw��h>��NH��h0�.� M�Dת��s;�������w�^��Py�w7�Ļ�q#�\�}�`�ZTj����]b�<�e���)ʂ�f@���F�C�� �8��Q�1����g	���/�p�����B]h#�d��N���D�g�@C4�Ө&�ż���_6w���ì��M����{x�f���HzS̉F��pV��e�ݬ�L�>d��i���92��.�
��_��·����w^<7!��m8�,�љ���2�%Vj ���j�"���`wS���񱊭�XN
��n��q�1�}�$�^)Ӊj�e�̌o�Ǭ�:�σ��s)g1�\����G����1C��$_� ��@"������V�k�-��yw�?Y�WX8R~�[=�R955Q5�ng�(,��,51/��a]yJ�������x���[�
P�/Ckk���=�����5��!�P�C�Hh�3�GT�Xg��ܹ�iH9YD ��O��h��)Ak4����03k��N�:�)�����޻�F
�N���?���t���>ԶT��*���ᓥ�������y݃}nU�*Z���p��n��>��0"�	O�,Q=��mh5���k��J� ��[.�}��5 ��lCT�[.-/F��a��3��$�#Z�Qdms�Ҁ$]Tw���9^ȷ
F�e�5)>�D��^�;���<D�<���@��>�>V�̭���i�fJja/�l�� �8��z5�.�x��^�B��tF.����Hds�3�ψ���Ew>r�B�~�9�g��̐S����A5�[3@N�8��A�ۏ�X�����s;�F�ٔ�!�Hcxl������@����fa�}�G��i�����m��\O[u��C����n��}��x-�@�ڶ��{�<��~	n
�2{�$�=�6v��!Q�^�*mH��5uv�1C)�Zm�fS����4�ohGE�f/�$,Ϊ�x��pt�SkoF�o]E%���	�>� �i/DH^�����D,Vޫ>���%Ti�L�+d����ђL4�L�Q�(~>*�uu��P���~���� c$7%�9��1�D���h�}o�^�yS���5��Y"�����j�gJ�����c���CUR�tH�E4��U����-*D/&roԖ�r����zF�z(�{��:�+��r�������!��fe�A:�� pA���O�*9>s��{���ІـN�W�s�8���[��~"xe���d�L�N�$��cxHj�\K"V���f��0�з&/ؚ4�x�!��k3�PV��nvmY�jJ���N5$[�ãU~��w��X�H>���(��`j�ؘb�rl-���t�}s�����l4N�N���L�\�ϝ�C|��1�#�#������gQ����`=�~��-���p,c{E2����8X0S@U �lht�b[�	�H'�J��8b�\Y�-�e�r���{���opM�++׀�'B��5��<�N��L�۟NG�͊��o0&.�:��D�cJ��F�����PS����+������?�|ִ?�\lV�K�#8g)���X��eT��U�l�ӋcK\��`$���<�4��қn� �Rm>P���
/�V���$�Il�YS<�^�-ea�㨽�Udڗ��'�y��K�w�|$5ͣ����q�)(�p.]���J���z]o��xpZ��"Bc��R�^�	�}�7�8��a�ۃٝr�~�3�gU�Q�,_`�`�4�����9H'���j&1o8K��˺Y���Gtf�����F�4m7���k�d���?1y0']��o�����΄pn@X?��Y��X�|R�Sm}���3 W�)G�x_�EX���`�Y�-�D�D���;�e����GUS�^��9%m���!�s��\�A�FoW�?P)��]�lxaѫG��ig����ڨ�B%���\�g�3!��-�0������� C���],��:�}�#��E�G�u��uQq���.�����Q��z�T����	��ҏ;B���^CO�����yT�S�:5`Y�+�d�T�q�39�r_��z�OD2������	��,hp�#��TJD��1BPs�	%���&-nm�>	+R$�Z�ZS���ϰ�߬}7���>%y��w�?���41|QC2����m�|^d=���� b"��گ������r��������������1gH��? �%:a
�9i��e5-ݧr>�)(��7S7�oS~�&��Q�����B��{;��B�A�����t�2��j����Tx	!s�#�θ`�O���!�Ӿ\/��X����V�5�Q=]-5��E  wI$zS�Q�_��I��;^"�ge�y�
�AL�[{b᝴=A�u�M��"��4W@kII�<��P�+�R�yoޅh�� ~�)H��gu��Uo����ߦ��Jn�PܗW��#uY��/�qPG?(=�\S�,�{��MiF���`N̼U�Y�mȘAb�x�Q�� u��9-&!�y;���O�}�~�s��T��͂�!��ym��g��8a\����T�VKS��I�d��>X�_� ����~i�9ŧ&؏[XE�%���1h��}�kz���v_�*E~���7�m��4c�C���i�K%D�� �ʽ���MkjE1P�����f������C������B���0=}Us5j�:��I��w�-����O��KK]m�2z+ȋ��| ���3�76�w�w��Z�+연��d���9��+{�*�o���ॕ��1������hD�Դ�>�6{.�0����t�܋���H&y��-D�%^G��,�!e���p:�F�����E���Y=�)���y��;"�����(�W�3�	50r����L}�҅������TE�,T1F�28D�I΢�qCR���A"���F]!����oh��dkLṣ�� �y-�i@���^��I��0Wo�a"v���t{� '�k˻N&��2�ȅ>od����:4��α�q�a�RR��\�>���{R�'�����Jу���؛u�g�sY�[����֠��r�������U)���n��p��������5��I�g%+�ټ�U�d�5����-�(��������3�ڱ�i�.���"(`���G~TQ`�͑���;;Z=�Y�A�e����2���Z�d�����Iu�ys@�ﱁ��L�ݐ�>Ʈ9�!��i>~�)&`�6�1/�J
��#`	x����`�ˋ'QS ��z���&7�­���B����&�1�i���T0�m�����O����WR_��7G���	%E�S?W����3�ZT�쎄;׭;�<�=�h"oxtc�^�6�����B�5FWQ���+s��RjL%�I��4r6;��4�¯7-ҽ&3�%B�1��c���G2-¼�Z��7�.EYȍBklXY��%��dx�o�x�U�#�Q�}T��E�2�p�E�t����͎�
]M�O䯘�B�:)Pfb�҅B��cNɳ7}ޝn�*�����+��[~��\��=r�py���Q�U���e��NH � $̀�h�v���%��%�g��1��˭Z�Y��/���t$�e)�0ͣ�7�� ASA-A�h���b�Ю�[.�4�QԄ��0?3DÞɭ�*���x�o�sX,1!$H-�����'.�v:�y���g<e��D/eͩ��F|E0�};?}˶4��?~��O;��6eܱ"ѣ(�B&�e\�/_VWN�����]{NS���5�M�=�y(��9��zO�k�Ps�\$�sXhe��Ǎ��pe!<�y*�KѸqi���C�!�����=�XE��Da�VJ�]��%��w�C��~G��v�^��*�\j7�7=I�+P!w���nB�	�Y�����#��7�p�zkc@��z�i��U<O�c*�����U�y(�:=� �&\X���y�ʕ�w���y�Vװ�e�[#�\��X�AE{�1���Q�q�����Z�3@L`��!�.���3A���9��Kx�Xe����ή��"�~k�m�Y��1EץXڴǿ�	'Xأ�Q|������sLd<%���c����<Γ���7�� ٛ���ϲk��p���!�Ҩ�y�ң<�u�0C4B*����i�L�ӎv��b��&H��U=ql%�7Jv�B7L���DwI�*�M����`�h\��,��P|l����,{���n&�|� �?m�K]�n7R6���l�Z+O�O�w���o�k�I��V����u�wQJ1����2xŔ$����U��~"�9���#�h&_=v;����(�.d��srtI5}�nB��d�'�T0B�̼$��%��N�4V�!�g��4�p��aB�*s���n]t��f�IT��`�@	�V���u��_�T�;��\�.���/s�n&p��^��"��!@��3A5��>�K�M�	���vF��y����vV?F�kQh��pد���A��2�]r�j!������	2|����$h22��Li�h�-���ۣ�N}c��K=0V�����P��?h{X
 .4��sD�ؑ�G�@��Z-@��}����Z郛�l%����3����T����гJi�ۤ �S*�H�(�O'�c�k��Ֆ�޼��M<�"�ژ�hu�Z�b�j&ͭ����#���v�u<e��517�$���ŏ�`�d2.��������e̻�>�ɸh�@�6]���_���2Z˳z��4�(�R�mt��3�#;�׬������䊃M<��ߔ�&FB1>�帊��POv:��&q�2� @Vw�n�A�^���@bx�`���詸�S��� ��`яڽ�yС�wHϢ�!��K��k�ٙ��;�m��C��F�/�~J���7�q�H�fjΡN`�ji����`��mj��.IH����2qV}.�o�>��+"��x�OR�[�����z��˗�<2o��q�UД;�@ǈ2wr����g]�v嚕� X�,��f@���Y#�&b�+V���͹��������c���E�JV��3�6p����{FE�-4q�*�>Bs%�+l�i��݋E�O��U*�����F�l��hI����E��m�\� zd�JX���@j).V����z[��hEAE��W�����D�V���&��:��9�K���A�JF�*�����P2-S�v�H2R��Fp��{C3�u�f{hroȈ����H�N!�d�x;��MVWm�o��x�2�=���b�4ǅ�<+�`w�n���z�~�+UZ��kK��?��н�G�І'�8u���H��4�D� Ç����V,�3��wr�W��Ҳ|�ʸ���
������FX�J�:�)��l쇉��\U���:pߪ^���h�Tqk�`�wi�J�Y�l�s&O�O�#eP�YL�{�r����B�W�|���_�H�=��~�<V��@`�*E����b�� ���l^��'�Z�>3�Q�Z��A�-��?����Y�}+��=��`6���1�D�3h���I��#�+�U��W��؝��g-����������"���D�A�q�����>��W��ȸ��n4󄰔��L�{8��Xv�%������p�:���7��%�)^�)^�K�1��*2��E�$�%�?J�É����X,K�Lܪd���)����XߴOu�)�T�\,]��؇�����m�*
��,`�w�/�A�T�Ip��3��J���Tt����8�d ���!�=�Ѓ���"R��%�#r��l"/��C���
a�Ⱦ;�^<���j+]�Ր���MD�x*̩�f�o�����m��@��^�eBW��YL�n�ri�J\43�(�=}Q�C��_Y	/2y?��SF�~2�hVx�2��j"Ěcw���\Be�#�عv��w:^���\	ǐ�9뺢:3m��FΣ��PU�z���EE��.y�����������5��R���E�
yp�\]�)�,h`Z��XA�-
;���эIir&�J����i`1r� �ݰ"�N �����]�N����n�%�Cwm���h���B���M,[@r�*tT���Ջn^$O���.b�H^�}�=D9)��o��:O����rN��ۏ٩\����Hၯ�/��w/V��8���l�.2	Z�f{J�z�y%��c�(�ZͲ�f�Y���v�D�ʺ۪X�	�LKn�A~��"L!�E�Q�5�-��#4�^�U�(N�Ij.?�U�o��	�3�~�ǥ�)��	*H�X��W�KGh���7`�����El�����k��
9�|�@�f;���T��'��;?ė�}�w�m��_��f(��nF�O\���������|ؔ$�mԾ�!�<��l���'����_��r}/�#���}-5Ff~�n�A�[�X^e�S�5f�}��RQ�?t!q�Q`��U�i)4�U0:��1}v�$��k���IZ�7E���z)0��QF)��������)5��et��_�d���0�O�.�t�����h�߄3�����}���Iz���b��l[7e҅ʢJp����>�kÍ��E�[E�l4FTh�%�~Z(�%��4�T,�� ����%I�.��!>�D�4I8�����+Z����l��[����A�à�7��ٯ;�R�>�i.hc�lr����O�_�7��g�p����߼��@�7�7���.�!Ւ��,�&y$ˬ�x���lSa$����ѪS�����FP׮Q\ί+������,������D\G�J׫-�d�1fLX�+C,<�&���^2Jv��C%�^��~�y�����&w���<m�աm g�+�;HE�`2,�\�s�[f����ց%��y�п�Ӎɺ+x&p�PgIQN�1ˠ�U`����Ðt�"PU	��R*�FD�q���jǿ8�yjz�V-���w*'^�o �!ٞ�h��%����q"e��A�"�S/�%m��h���?��+#��[��z2���
P��pٮ�R�K��vb�Kg}�ó<�1��eҋӔm`nK-=r��SfI��g)��q�iH WZ��ȇ�hkڥ��ҪPt���\Z��:�fX�4�}z`=��3`78���(���̔WZJ�n��u�X1Ya�IU����8��b��H��3�;��V�}�b�w��t��)�^�Ȑ+Xeu�|H��+q5q�
]MnY�F.n��{4ڮ�!������`���i�%��|�*�GB��	@��:n:Sh��rHv�a��*LF`�ayh猢��0�-,!A��}|Z_h���}�%��T�t���m��G�%�ڜ$�X?��ަ3�Ul��n%�	�BsE�9���������m3^g���/u�&�W�;5c���#�� �)�����W�s�Ϡ�y�.T�tӉ��x��
�#E����	�4:�H+�W�k�F�q|�h)���ꢥ4(|+��'M2J�";��~��13��`.��haSs�,,����}N�e�~�{��V#��;-SK2�^�V��R�IgqʣK�����7ŷ_�'j"~��]�R,I�ç���P�whF��_id��׎��������9o�-ſY�	��xɡ����r�H��|Zm5� .�"�2�G'�`z<�ur��&��U����-'���?�!;����;��X��������ߔ)[1�u�>Y��謋Չ��Y�"���:1+�$��r�1������3���}�Bse��(�!�%��;��~������}���}���_�TRK_����
���2}��
���W��="c����x��9'����E�m��9��C��U��t� ���.���KԢ���,���w��D������������]�Ff�XA�ⶍqs�"ј���)�i�-���/�Dt�)�Ė�~�@��t˙y*��A'0-,�3 ��c���I��$�P�8O��(��"��r���tR��d3�uȕ��?�������s��N���c���$؏
��d�`�ؐ+���K�8)��~#)#矂��'��Q#	o^E��EL��GޗiwG|Q�l���ΟSls�����e�3g�!��R������2tcHL��~�����y��u�O�}>Gܖ�p�$T@��q[�2��Cr>�=���æ�`�Z��T���z��Ka������)z���QQ��B��.$�ً�u�n��6r��0ؕ6�+�m�	~㯀�[���ě����
"
��$�%WN�%�iE��hlMf���jґ���� ���@妇�����1�n��2�p�*5��g'O�"���y�ɫɜ2#{	�g�G�r���4D�>�1k���6���P�n�H�<���u����Җ�/j&Ox���p�.u�30?��`�6X��TN�r9ճZ�Vg<%}hN#�J��Ud�I���O@2��]y��U	Eŏ�9���d��>e�8i0�gmr�g��3��m$�_#��w���k'���٦�K����o�NR� �����~�x�p�rH}ڽ{�\��B��u�d��O��/tf�6�(�O�Vu��%�*FfI��L���l�����U/��i@�a�o�7��j!���Y���ϩ�P�:�8կКi3�����d!�[�Vϵs����2�����R�s��c/kVzT1~�"̬D,xM�	�$U�Y�r�>Q�����AR��~��������q&c?��e ���L��%��%�]���������c�=�iJq��qX�	��gy��r�R�7�'	:5I�������&�c~ |x���s���G|{̲�?�3�}�D͠�~1��P�ܱ
`�Myw<�z�n#i�d7����tHք�c�ᶟK��VK�@A����C�ۺZp�D��c����8�L��?��b?d-�D�3tg�Կ=��f��Y�+���BN���Lx���
Z
�/w�G�מG���<1k���%���q�����㗤�n��r�h�]�sa�lR�b�@`����4�~H��!���KͰ ��gECi����Ǽ�	��)�^q�G��lT6�0sf�3l��&l�B
�p՛G�с���$>,�	�5�4�J)q�R~�7�*�ב��(�e����7^�7|!�!E;	|��Y<$��~�'p�@��=�F���Ԓſf��H�d���k��-��%g�͊���4���ʇI�Eҙ�����{d�������۱���.�_#t�r�\(�U.�1s���WT���e���%��	����� ����˯�>R�d$�0ҷ|���n�r;�)y�6M�}������|=��Zm�
T��*�c	B`)�S�=��)3ANv$	_�8���~�eC<��&5�\��)�s��������i�L�C4α�U����`J��]�Z�`V��}H�6ڞ�k�fU���-�� �huJz�f}D�R���祐
��㿾���f>�wi��y���'�*�/�K�S��B�䩐0t�TV,w�/��*�T�Y�$xf�R$t�/��~��@H츐�C����(�ˀ�E���K�Jq�;z���������H��Rܚ�q�NB%^���r��.E��ɢcqf��A`�
��~G�'WG+�kQ�i!�̦}��H�?e+�A��嵎3�,�bwd^i�}G�Z�y�vtN��#� � �I�_�H5/g5Mu_�h?C�s{L	T�B����Tپ����#b�j�t�L.kw��{�|;��Lb &��q��U�\�G��C���+r��)U��F\�L �̪|�\��?#v�(�3���S��8����`��Q/N	`	y���(^YU�Ŝm��Z	MPvTઔܮ1��gܔKR�NS��d vP����1�܂P6⎞�������㪽1�{!&ݒ�w��x[���K߈\��8�ɗ#z��`�_[*L�����6�x>�9HE+��0��Ws�F���H�E��Sј:s~���3�P:�����3by�_��֪vS���y�w��ɥU��ׅ�e�� ݍ᯵�ɣ>���^�	��2R�щ��۞M�Sԧ�+��gR*;(�*�9G�}ff�H���a��$*Gp�(����'��	5ے�<o[��Z��w,>�>����L���4���*����՞��!�!�<�Znn��R����Z���w�+�}�P���- ��}����sH��6�3�kx������hMT6"�]�����3Bƺ��y=�=�l���1�) ����v��}-#k�����D��Fw�ko"���-:���½����Q�s��V�;�(�m�A�)/,-h�X��V��$lm���kn8Yb��%�
|�My3�M힝~oe1��Jtd-�G���e\��E^��Z�-D��l$v���<�pι�a�;�}��e�gc�Ŀ55��k�|�M|����˗[2�����12�ߦ�ס��\�{XE���d���i;�(�Pnl�k~��O�+&{�(�A�uhAt�*����t����vjdi��}��f\�k� 2�C��:8RI�e��{���nF��B���E�<8����K�b��oZ[��<�-<��� �$~z꭛�����kc1��Y���`��K���o�"����@䯉�o������Nx��y�<�Cւ.=O��9	яDg���K�d�������i�v�QW���nΌH؄ڗ6&���e a�!Lϒ�kϥa�i�ZBМ�^j�֥^��4Ol�^�%��]���/�h�ݏ��て_oi�_���:�G5����=� U��@�Z��������3h�b4��I�#�u��*)ųF���bt���"d6�2<��w�`swv#���Nyb)U�Y&�H��!���4�ԻrԷQNU�Q��+�$H�x�!hｊ�g�� �QzV)9/��\s��<��c&f��h�w�]$h�����m�UM�����%r͔!F9ُ�T�˂5/A4w��IdpKg�=}�\w�_��Ou� �5o�CY1aTE�ڽ���}6��5f	�9�Q8;�r��Z�&/��� ��|��P�9�;Y�߲?wͻ����9��~�i�t��<�*?l��3�y4.W�`��ڛ9�>;��������f�q*����<_��z�J��d��'X���#���������HW"����#����� p}�K�,>��+u����Ղ R.��̎�w@�㏕p��{`�"y�f�da�N�A�쾵�|Ƅ���N�au���9�ҼVq�t#�������W�:S�1ۦ*c�Y���:^`Mz�6lG�]�a��<A�x���mVw	H��K�`Pާ�b`S������
=[XU��EE���vV4���Z�
��ҙ���wEw��)u$�`xc���G�Ԟt	?ixz�D�@js�rf��Q�u:���`��\��&N����@e���p�5ψ�.4_n8T����)�I�T�C�����~��$�|��1s/����F<��{^�Ӈ�@Y�T\_^E��T�R�?��
,�}�d����ڔ�D��F�:�g}z�;�U�~��h�e�R���#)w�O�,��#���ԛNa���)��E��{��i�\P7:�")X�is 3��w$&IZ�k2~º����9Qp�9�:<�Ʈ�Z��
3�_�
�L8��m�~4!� R�Λq>*C��X�P#��E"�á��Ħ=z8+h$<�z�z[ZA��0��}��'��7�ot�?w��B�N���<��<�F�֒2��	������1j��%LaC�k��O#�YB/o2>h���:Ƶ/URQ�n=�����X�c�k��M��Ch[��� l��~i��?�đ�I_��Oƻ������l��YD���s�^��j�4�4M.��N�3���o1�Ɵ����e�� �c�e��@g�a-
T|?�?/i\�+�A�
�\}��aK�!�>y53�I~���O�)=�^����,��H1�-Z��ژ��"�X��p��)�+�O�(ܝ|RQ��O��**���2`�@$^�*��+Y�\��^= uD���	ck��+�1Di��g3�M u�8߾���T�
��.bɼd��"+Br5x
1*����,�rg�
�Ϗ3�����^��)�^̠k�X%b|l�ܑQG����ƛj���;����nj-��yYd}�ҵ�J�D`o:���]�K�������l1��Ɓ�ˋ���Q%�M���m̥�Q#�B.s�L��l����W=���
8�D	�O��N��~XZ�z�{�����
�������b���W�雴��-�
��5^�
�B!����'��'�-OI']wߨSPql�	``�/�V6� ��DW/�����I�O�}�q�
^T���2oaqo!'���t��-Ж��T��8��&�m;9� �U�iͤ"7c���萎M�֍ø6l�s=�I4�b:7�6��y9S|Mx}
�8r,�F[rHoEU�m�j��ҟO&7�:�������G�&T�*/;k�9��Jr�$n�)� ���$.��3}��o���έ�����!��MH6�^�"����t�[�-�=�拪�v�CK"9��욊 _��rva���"� �I�w��� )�'��u�É������C���
D)L�(}x����]/q$j�TЁ=%O��u��UED4�3^ȷq�����ZK�jl�8���;d�!�҇�9����c+�P����$�Fc�	� ��
7y��1XQ(.F>dA�����:��6C�C�uUޏ>�&$p�9(
���I+�IKL�Ȅ����2�� H�U=�N ��s��m���FD$�xx������ ���?8��z ��Sg%�,�xY��2�i*s:���m2���9|�yn(�#��b&�쪏A2�&�R%`pZ{$�%�ā�B�t�|M'�x�ZG���FI��I\����w �3���l����^F�T�U�H�AoH�2k�Уr��HAS^����w�$�R�J!���O��!v��v��4���N�o�8<��(�P��ξ �@��8�+c]n]u�[I�h,FZ����N�B4[�ģR���6�����
��/��Qn��_�{R=o�}�<dA8q�O��Ϋ~;ٶAlj�$]�u�-T/
j
�������<�V������P.'?�*����@���yd�У#��i�8�+M���7-v����9�K�*א�����\��o�1�z��´a�NB�I��wҢ������<A3F�rM��t�E��e	��T�rC\B('J��촋��+�AfPI5O�a�ȶ�ń�}Nz�Ã�{�s5!�x�t{����Q^A�~�����$o���]K�t���&�r�tW�I��O�!8�Г���'��Gټۣ�ۊ{�/m�,��È���HJ�Nȶ(U��~x�x��6p�Wr`
8��Ion$�8d�ա��T�K%YP�I8�Z�?��@S\���[}�f1	��Z����:y*���roQ�D	3������O �l��I;�|ko�1E��Vv9��=�`z�����]�m��>���.�y���U��x�ÝmZ��3��"��7-����5�]��#�uf�䛔�0�,�2���M('�',�?�M/?&Wj�Hן��YN���m�,m��:��A���gI��;qb��?�����?+��ⱶ�g=�`�������ɽ>x8#����zӋ٭��XiL_D�7�9Z�t����l]u�hz�(�[��?c1
�w�;�bCR2��Sz��Ģ��p�֋�S3���ȍ�݄u�"2[���I���}q�p9�T#<
쌳S?*�
�=��w�w�>�2�L!V��A�Y�Gq>ܭ�Ŧ;Q H�fU�5O�;�lR�1�Z����LTx��7�R�ݥ����y�:cB�H�n��?H�tӟE1���������F�.�|�)r1�H�ι�>��Ԍ�cP$�b���5�w�&���f��s5C�^���I��H�D캡r� 1�/��\M�ڭ(���Zt��(U���-��`**��D���6_׌��U�UL![�oO�*_������mB���RJ�.]�¿�*�\�QAC��޵�;u�y��AˑOׂ�^���M3@y�ێ4�����&�A#]W���X��MOv=T� �}\�ρ6���5�������Ýʋ�u���D�N��ݫ����џFôlN�29���<)=��ӣ`������<��Ԓ�~MM� U�R�F���m� 
t��v~��O�C{^# |G0l9C,�kd9t���oyTڨ��$�fԑ'b����G �,�=�	��١��.2/��6i���%�]��bK$��+l�9�7� 	i���W(�,��9�^0�M����4�W�k�4�$���Z,[9�S2���+5�5u8�(�Q����H��0�;O�?$g&:��f+���Mt��7��1���"��*`R��5l[��A���P1���N����	vO�gm�Yy �-6A�!MŷD��kQ�d�ꠂ�%v!4k�K�4\pBOT|dR�~#mC�]-��d?C�<i�'E���U��G�_��͉�i/Q0��#�w�ÞLQ��ލ��,�	}��=40ϗ.�ٮ����7-�O�A'�?�m�ع���^���KZ�����,�,��FE�d�/�T��xv
��5��#'']&�RO�F�*��m਴n�(B9?�d>@pEPV�v���x%�]�6t��﬩�c���Y}�g?h.2�t~v���Vn"+N����U O]����17@��q��.���C�k[��%�I����VV7�	��g�{'�$&���4�5;�|�*Zs9-��'���G�� &��}8%��j����D�":d��"�sf�[�Sg<�xqj늻�:h.M���P�*���1u�؝Ŧ�g����@�~|t^��G����A�f3�,���m��)O���ɴ�C�o�-#�3;P>0���ΐ
=���a�rh���^f��ӄ�	b`u�e9l��ǿG�q*�;�l�A��$�g���@���= *��f�gR��z&+�}���B���]D�:�a5[7����|����Y�D������>瘾����h9��H@_�]Â@k��av����~��q����ǖ����1?z� 4e�S�6�R�dv�v U�Kؑ����}�XP�|UIm�є�~���X���Զ+H5�f��se�Uq��q�tD��d�}Sw��{�dEõF�@�{4ٞ��3>d�@��P���n��2�����N���y��Y<�r��ٷ�g�L��� {;�&F��P7/.D9�>֣ �,W���1�Xpթnb,�Q~l�����tN��t�b��]j����_rv�uT�N�ٱ��8z��B��c�Q�V�ɆͶ���b|G|�j����3��R9�L�t�̻(ȭP�%F��p��#���v6�^g��\�t�`�,\��;�)RP,�[K����q�����p�� ������$+�z�-&��#|�.�%����/�'��$�4��)JS�)�$Ĭt�;j!��. �&�¯�,�X�m��1
�ݞ�a���ج�~56��r�緞�h=+Me��TgAڧ�#I��6�����?䓓w�s��A�S�x�h ��<�A�a�����\��m�"+Z�s0=�j��?\�P�݃�A��n߭=��;��{i���a�m�X2��	�󽵪�i��c�+n(<��'	��o���o�>1B��Z1�����y���踂0'/�Tc���u#��*�DFu`>�U9�O������ջ&�U7	g���~�� �,o�� ����1#��P:�\����&�����Ǫ%�`����8�K}Pwe-����pJ`?]G�T�(��i�:x�qU��N�&pIr�m�Ф���!�hVe��0Q�B���g��Bm Sp��3����cp;P!�?��s�IX�	b�5�gb�T�:❍X�oO���S)�/ �Y����bwI���� � �"ֽq�ᐫ2R#��Y�Y�X"���k� bdV�����S��i��%��w��k@��Y��M�\��hs�0�/�Fz�| [�X��
ڞ�~�3oe��FUd�F���c������"s�pɵ���-��A�%$���`���Ju ֟�B/ĜJ�)�@��7�R=(�hB�\)��%��`�w]\�闈�����kftu(�	f��0r6��\9
��9�s8Ր�֣��k����R�����ϷE'���������(�S��� vJ5�;�-h� �<��� ��Z)��ڢrO�
.������˜�Xt	b�1�K.���x�_M=6I���"Ҍ�+֡�8�2�X��n���P��ģF�6�y�n�s5҇�Dڲ�&���a,q�:�t�˥����8IgH�Pذv2�zf�����#��
��Hj���i�n?`_4l����)!"n~��)�gʠ�x-Ɍ�J�x��-L��v�]�j��5��� �L;@��g@�iͫ(�8΅!B�ʳBR�Ղ��0�gۘԤ$��}��V"�a�G��/�l~6Q�D����}ࡩO>>��{���rާ���q}��H�������I"���ʋ�����~b::D�j�[���Wd��%�[7��&~�0Q�u�#]t�L�;MeP�Y*U��Q3ma���Z�����<���9��L?��"-B<�xd9�x�p����=G������
����~3��N�+����{5�v�m'�����1G&x� ��z����t���@!��sj���(S�؂���6��(>���|��K�&\	�NP[��n�t��N�MZ�[�X��q�$�P\�:jY�.�2�Ȯ��Ye������v�
*^(5l!����]��IsEg0Y>���ᮇu���5TM�]����K���,7�{5VP���iPA(��~����dY!h$su��psE�jr�K�a�0�_����1�t��]��Ļ�v�L���I��R�M����Y�M�4�?���߶Tx�\����/���*k�������&������ �@ܺ��������P��-��+�j6Ly5mE߽�Ԯ�h�x������x�*e�u�̏mR%>僉���*s�u-�jk:����.��#��K��X��H.m(��`g�(�y��3*���jh����Ey}��>Pq��$.5H�f����������F6�؇Y;u���wh��|.
^*��*&�i�L�|8�d:ћ{���K�2,���	/>D {`,�����-�a�`�g���lS9S��D�4#�_�t��0Q�-������ԌX�����gX��${U���)��kdS&(�<ÂKP+��%>��K��1����l��Ɛ���~��o��,uB�޳oT"� j9۵�q~��2H��U�G��q���u�E"�;�N���w�!�q�g[8���_a"y�尯��u]��S�s��i�F����,�dc��]�H�N�5PQ� C=����ϭ���Ө@��yvflr���$�b�"�d���<�CW*��7=�htH��A��M��d��nC�g���~�}Pusm��R��or�<HoU�j��q�tp���j���e��^�v��j�!.��3*���q���=\�]�c	�E�B��fiJ��РWc��@��˖�e���/�s!�Yx�"D�h�h�.�U���e9�23N�2y��:����P��a���Q�gFr�>�}c�I��.���6pr;�&��K(Ry��m,2b�ؒ��g���΢������mG������3��0ܮƑŌ��pRc�^����t�9���*��g,_t���5o& �ꭅ��;V�?����c������G�3(�/jA�d�&�{�B�e�-{�W@�gBxHB�8������x�F��y�m�0T#�?{�I	2�v�]�w)g�-��C��LۺEBϏ	�{�jo:�� �f�k?l���
$�Ĝ�XS��}o��_�)뮃WZ�)���6�~��ݪ%��(�:���7pjur���l��
=�I5d`��wˁ�� v\�����Uj��3Q���`�P݀pi�ْ�ED�.j������bFLQ�q��}���HM���e�U�*�lV;	���?J"*f>{1:h�FsRA�ݠ��d�ٝ@�8��:�%�M�����90�hD�o�!��pn$Y��]�s?��}u���u1���qn�9�i�v)�G��^�I���=\��ցO"�>��%�Ɨ� @a�u�X�{)1��%����.wq��v0��v�{t�����n��y� ���6�:��J��7�|�1�8�غ:ψ�dbf�+Gs�.>�+��Tpݍ���F�mG��c['�T2���X�܄ҟ6�O��x|fР{%�s����ᴻ�Ŭ�}Ĭ~@�r
KN��]�Va�nX�G�V=���]�m�8o�_��C�4�K��@�J���H�� ���7���%FAE`�/	�pV���lG@}���վ��R�\u!|>Зj_2���^+b�W��z ����5$�*���&��7�h��S�)�8�a���VC��I�[�`�a��|�����{G�9�2�9�/^�p&��Kl��(񂪸8X�x��"!�8�/��aS7��K�f��Ú��a���f^�Oz�FOD��Ӝ;j�����Q�����7���6�}�q�L�DVH�a������*�{��ؗ�)A�su���s���=��KWӥz�(�	ϳ�,�@�6��<��C�����u�o	!a/`,ұ��1ա"��*��t{���� ���Ŋ���9�rG�5�S����N,+���|�,!�&�/�f��C�I�,�pҾI$��X�T��ϳ&ܦ���eO`E'9������ �E\X�r����~�HkD�"N�4`a� v�k�&�Ƌ�&#�(�����TS�5����V����Jtf){�-�<0��H���:�������u~�)�(�X~�Qc�- '
QL 6�HH}��4�X����L�"@@)��1��kU@�j �����\�i��e��$Ǽǘ�>eq�?Y��|1�2��,%��0cq6U�b�I��S��_N 55'P���/Ѳ$��q�5��E��-��k�������V��<���Q[<�Be];���j��s�FOmPxұq<�%�k�lb�H:�߮�8�a��W��nמQF��M,E*�"��"v�9wl���BƄ	��� ����1я���?q V�<}��m��<o�a#:����	��	�G�!��/9�X��m��'��@�����Hoy�ݒ�:N3|nӄ�����<N����e�0� G.�z����%n��n�`&�^6�v��w��vD�3BW��U%��0��%-ݳ��zu�Gm���㼛�Q�5$8�K�ʴiX���J8fʍ����w�3]y�+���b�-�^R	I�>��jG�h�N"��Ϯ���x��b�ѡOK� ������eO7���3A*~����Jݦ�U3���b���-K[������`��������:��A��&b�A�%'��X��f'E��1bSK�mH�YR�vH�=�S�:��|B�v��ft����#���i�%��^�K�N��8`�"=A�y���f�>B�tTf����JǏ\:q���vS�����������\J�<�vW���^���u&�uo�折�EE����)񆧆S�k�B�tʜ�˱�y�Ǜ(��Hz�^��ا��_@w+7T?)��xg"5u٫���o��rO.�L7nLN���:S��Ӻp����Ԭs�$�X�㽒��.�����-��w�r��住�g�g��)/6�6��\%w�i�Y���:93��t���@�ĪJpG}[���~�8�)���\Lf��U�1���^�)4�A�8�e{��SLK��>�b���22"01H.���t59��)Q�����{�e�9�1ߢG�)2 ��
"���[Iw,i�$�i���} 8&��u���	a�FL%�v�FM�E�N�Xm����4c��K	u�̃bލ�br���C~�%h�>��)��ݍ���6���.�uK��ZE87�P7�X�"�a���d,[0�2H����1ݝJ׹ĥs)��DF�����j4~�xv�0R5�W�����חj�D���gHf���S�uf��T+�r�<�]ԭLG�<��@f/��I��3�_�5��Tf�2���DkX��~��N9yG�����'b  zqit�p?H(p��5�����A�@��-���9�cÐ�Z(�p"T����f�@��&\i�����R����.���{��!؜'Ǵy��#�
,J߮�r
�ǿ����$ ���ǚ�7���Bϰ���?tکЗ�s�����$b�g�&�M��-#A�[!�� ����k�m(R��2�,�䙯B߭���\;����NN���<hO���/άw��1�km4y�񄆢�A�XŔ8��x�*�������[����c��Ϛ�[:hys�ev)3��tB���,FtA|2�\�[,�@�"]��9�n��e�ON�\�Egaя�> �CnF�>�<Ȁ���`
�Kž#.�i �����>�k��C��}+:������&_)r�s-΋���ᬰ�*��O�.�j���i�B�j;��Ǿ�/��J�e�-�ۿ�,���2B�� ˱��c��~�û_q�#�Rfh%I�S���������7< ����_�Xeq}w���C�*9`*���c_�"�}����k�wⓨ�f~���)u Io'�L51�t���%d&�_�7��N�i"���*Y������ &F$`�¯��8�[��:�����-��e �˾_���:Ć�����K�ҚI�i���ua,�+�u��S�Vd �c+�$��H�:�K��5q �N98(�/ӵooj�g(>���d�/�؉�'�ItϢ�߭d GI2�D=Z�T-���������6�b�W+�T�/l��m��%�'�UEn`����(��BW�k�(����s���BkK�v�0�{,~׏���;�����1E���>�������.���Q����bA��؇�<'$cŷ���J�-{>q��������x�x�-�V�7u`�wz��}���{z<yD���ߎ��\��DI�Dƒ�Ƣq��C��RDv��h��F	CL�w���8=�g����������)o�,�}�m�NH�՚�����Y�����\}=�����U,�ab��b�s<H��{㐖�v�C��=���!h���	�1]f�h!����gC�e���(}zG0pl��C��{!�Z� BT$��8�����u���/S@�������1�����qe�o�*��%fU*�l߷rv^15 ���=��9�&��\�η�*Ztf����T�0�������g��Y���4DK��-�-f�qnIh���(��*&CL�QF����7(ɨk�yb ������X�(~߱�O;��4�_q�a����W���92K�[u	�`Izl�IHk�b�H�OG֡Eu��*��	�+|j�f��e3T-���o�]F�#���rzo� l�.x�����i�K��)nzJ߰޿�F���lbN��r�
?]9�,�����Q,���H�#���~j4���xG�ux�o���P�&ď#�0u�������D}���y=` �bu�o9YS�(o�����e��� RwA` ~d���xG�W���X���`�f�^yN*N(gy�R^��6���7/@?�l3@�:ڥv�i݅Y���6Ţ"�n��~(5({���D<�b'�k�{�(��6�E�45:x��q:yTR=ˆ��Z7R�im�%ǫ_�_�ŉ��Pо��J��=�ǲ�] �z�U��	��]c��M9�=}͝����d<�T�9x���`��Y�3R�@=����,�6��G��U��oR�j�X-2r�]�9lfѝP=�?7&ri����1����$�Lxt�_��W�B~�Q�?ϱ(�?�����H�(�����q�eb���
��C_ӜUDؑE���~u��ͬC��l���7������4m=��޼���������c��Y��L/߰�܊�b�_�>�#��nݖ�Se2����W�t"Gzw���0���-i���?]�Ax����t,fEO�ؗ�ݬ{�(0���qe#LYUA�X؞�X��|�Hΰ�3�[�m3�lݦ�7�r�����Ť���fU�k�n��N,��Qo��Β�z�/B�3�<���e u𺕸p=�J|�Z@Hl�{���9:
J-L��+oR�0�v��A_�����@�z��0#���Z5cπ0��sAk���� ��G*��o=���m��d��ˌ3�"s�)��a��a�W4��f�I�D������_t76Y������J�����Mo��=�A�t��X�%��!�Q�H��b��Z�(�e6;��#L[o_�0Giu�c�K�Si��,��w~�x�� uK�l��[��.V�Fx�x�ȜU8��7z�<RH7{<������[�euƣ��@WN��\o�\c���F@�:vU��r���]Sc���8��d��${��Y�C8�X��ഭ��^��������y�f<p���B�c
N?����.SJ�����!�z�#�Y�=
B�(k�4�l�0�L�b�xZwi����4��TM����~ַ64� �N�@Q*q�[��Kڋ�.[�N�m�1כ/����I6�
p�ܝKFi��y_(��D�Yr9��Ԛ
��]�._0C= ��&���H���?�όWR��A�[����䔘uɏ�w\J4rPq��݊	44���3�D%/c�T��o�ޞh�U"�:"DY�f��
��s�������Uދ|��������U���)�����ԗB�I��~��_��/�X��]^�2�L��� ֌�G�L�Xn^��-��G��*	ɶt䥩@�S�@P9�lJ#�ٍmvi��*#fb�rV=� �g�����95T7A�v���~��2��4ߝ������޼��!��ZH�e��!%�����!�<��ib��y n����`����U�';NH6�j���ɧ���o�����_׫��J�����C���]�9h���:��Cf�G�.W� ��`���b7%�O���$X[G\�gc=(��/���͈�~
!w0𧞞�f&g�C�e�\=8̃���.	-Sդ�-��|7u���Z�a[�s"�t�J���,���zAzLZxf�*�l}��O��5$�S�+jnu�i�n��cz�����,z�,Ӹ,�U%���"�l��ASo�����퇩����y��G��Ē��9)��-ٽJ�r������vFWeA7�P%C��.G!AD�"լٞ8S4u4��=�~9b��PH�w!8,�Ő���\{�U<zQk�)���B�w�k/��Z?4���� ���^��4'Cm��|ƭv]�	)UH�J�H
aʛ�f)\��Ӭ��|!ē�A��[��E�B����sك�`3��Y�w�fZ�M�j1�����P��G� e����]�T�cY�x&q����2�^C߁�=��d\t�E�h�j�Տ��X�C�A2�/�?+tSV.�_��4�i��8���ZH+�E]�q|��5�m��B���}4���vK)�_�P��.��Jyk��}m���s��J��I`[�&8�^��0R�;�>�#8c���4?���3���)��դa�OK�G�W �!p�achd�B�!y�h�X���)$O}����ν%T��R��(�&P `^v�(r�o��q)t/��5��o:��E�\)y��*��'�ıǆ�d?�FD��
�ى�MbV��՞�.\>4���ȶ�!�p�{-Ig6N0 #O ~�+���	�엀�T0�I.�ɻZ�mw�A@����
9��l�sn#cZ���s�/"�8'��#�B�)	3W���<����RZ�B������bq��+���?N(U�������p�<�a>ܨ�KZ��<��Ca�,�1�<u�ދ2���ʵ�#z��q�/�ÓcQ��������� ��𼺘��'��0�o7>�@���Q�>���+8�I�\i�χ���G��t}�|�k$�؎s���?�����	YD �DM�?d�wꆳ���(=���D���H9F�gϫ�?��#�
�i�+a��e�y�&��D��'��lb7��S>�0%����7�nu ���bFL-�z���ٷ��.�i}-�?B�,P��mf�}���c�b�)��]_��Ǎ*�9��V�z%t�2��?,I���#�6kPiH�9~W=À�s������֤|�F���if�V�c�ԗ��x�6�y��Y�|y����}�C����)10�0�fY|�����/kV���˪�ϔd�hv���i�ț�`�;��s?[B1a@1�v����Q��[2vD�=�������z\5�X;m�Zp���H(�&�R�̘�})ZHU��+\�x���ЙP"��O][����4�?�m	��<c���%aTE���a�Y���mjrocw�z���J���/����7 �\�d,	sЎڋ�����+�A�/��,���Sc�$��T5ԉ[��T��<�+�S�,�yt�W�M���!����膬(�ݨF~�:*���w����{lTNϞV3NL��,>nа#O{�\���"�\I�g�ށ�m��dOׇ0���F�ѧk�� �Pw�9w`�M$/x��w\��Ls�]h�m<53-	�$�� �������X�Cv
[�U�$�qtvzn�
���/��B��#����Z0�u鸳[AE�r1�X5��a�3�]	vS�����*�������Žc���߷���-+I񗮦�P��L<�q�"v@\����w;l�dM9�\TF$���)�쟋�ʡ�������W�2K*N#1!s'��\��4��|���Қ�܄:)�/����aE3�n�Dx#"�|��=ڒ�;r����{��>Ps�C<vm@{�d�T�-/���h��}�[�q�2��h���+�h�6��r�oIu=Ph�m���8I�0�|����Ki!��Ka!2ή�>b2_qg�kzUZ�D�Q
O�������9�oϻ��X�hm�mn ���8�quH��G���fAggEת�@x���/0渋{2����FH�Dbm=�^�9fl�F�0?��@2��)�p��CLx�]����W��'�
%HX�_�)eV�i��G�"e�Y'D�ܸsW@�e�y�ϴ�����ܲ�T:Ed�AQ;<��RE���KPS��n{�zy��l�d���Ro@e
/ �X:���S�W��m���mx�tv$GSlώ���X�,�Yٌ�Dͤn��P[�A�^=emB�N�meF�L�-&L��N���؏�WLl��Me6M:͉����~0�|VB3��~<�L����+�� r�9�;;��|����6C�P��	������`��l���~b��kK��^s�qV�g�TK�Ӌ���ĵ���WQv�کw
��bZ�ٌv1�'#?�mϻ�.׉ix��;��B��y��h�NX�_��!����~��v�}ɪs�`U���Z+2���Kr��7 wL�5��(�S� R�]�����쵴�Nj=�BD5�-��o����gf�U�����
����؈�%}g�5�
�VD��?à��f�������K�Z�v$�d�1��_@�A���P6c��	�-aH�:�"*��.E�~�o�tf�[B����&t�6`�ŏ:\��صFeu]r���r��h��}�^��+�����<���a���zDN��u�ai;�Ș$u/,n�f�p�33���֩	)��Q�"�qb�b�k ����u�F�u-��5V贮Pl����k�W�zM��@��mR`Y�?=ɬ+Gp��#C���t�.�TL�5<B�X)�My��[fg!9��C�?'��P�����`��h�- ~7����8�qx{G�/�$H�jW�p��~��$cd�@��h{�	�P��C뽀7Z| bI���<�6��mm��x�٢a{"���iĸ��AZ�?ߛ�j3� h*9��G[�5�������x��kc���\�q@Jz�K0	��-0��fO
�Sq5�ͤ[�?R��R�x,��ˆ��`*�(�� a�g�@��Cf��"��C�~�SM5pSE�e�STj�?_N�Al�bO��R^MZ��nS3!�8�9� IS�"�n�^�'t�`��jYuYZ2�����pv7��WbmZ7��L9�	���"qu��\�RμG(����X�ˤ,�N/�#�n��(u��|Z>��~al�+	�.�OU^H����l��SFPE-�C��m_�m�cM0�[5��%��r(�]��m��T�?z�S��Hp��\@�K�ާ�#7g���A�~�y�f5���^�� "&aj�'v�B�)<��a�VB3eQ ���~쿿T�t��I]%Wͯ�g���c66@�B��{�Da�V �ہ�l��%,u�VH����r.4�`��z�����B%��M`\�.��� ο lI?9M���5wi���e=���Q%X��+gez%��3�>o��13�ٱ;դ�0��}H��N��q�߸�<���&kt��D!ǵ"����k
3�aؗ��%�k����Y��o0�'�>kem���_�/��\��i�Z�a$0S6���=󲃽��n��3(�'*}m/n�,��/�q�V]�J)��2y7'�_(`T�(�uM�jO0�&:�y���%=B8;{��%\�yo��*hwӐ����%��N�'���3aV�D������nSd)�2T��Y`E� ��H�稊bH�oUp�����5$R���\�y��Zjmd`�������`$w�Z�m���{BV�k4҃b<[�������$5�8D������,��,��.G<ۙ���p0Е���$Ƿ�»�oH硡'`cL�6�^dg�d��0�c��U0	ԥ���M�Cj�w�;�N�4�49w�U-v�z(H,��7|�"���W}����.8��<և.���!k@e�߫��vٱ���]Y�J��3����*���M͵��&g�8�N�]��7b���oT�.͛��u�~G�J���TV��I(�/됉��(U611���+� 2�l����5i�8haud5�un�uE��BQ�7'|����C̚�r&Bn�E{$��C%}s���8���̡��]a⵿p����R��5��Ѿ)#�����1Y��:�Aؒ�(C��f �F�N�������l���k;dwTp`\�O��F�R�.��Ww�d�mL�PۓE�H�F�R�<M���ׅ���:S-�DD5��aO�.0�����e""{��xU�L�9#Ғ��$Ȅ�����.+��٥���9��:���;���ic	�U�x�
�Ku�|AU�˟��B��M����]�R4�6��e���Y�2yA4򸢠̦������^+:�_�b��WBB�>+�d�������KEp�J����⪫�X�gq��|�p��؏*C��ZQwtn���b��� "3/#��z"�=|��w��3e���a\l�V�$��߂�:H��!��й8��2�:G[�ٝd�D^}t��#�Jds���e�kq�H+I�kn�T��_MH��6��x������iPG�[���Ƕ
���x�S�k	gן�3=�_��r�UE�Ng� ��f
��m��^�#& -��raV�;���<Nw7$zc�E��V�=r;3I8��[�n�0;SQ�߂��sǃh)E}_�S�AֶT~l���sM�?�,#@dSO����]i;{ˌ��p��_��y���˜�:4 ��r��Ӹ��3�:��[�Z��1)�p�!��޲�Z�l� V��3z���;��'?�䢚�h��*O��-g��4``׮"	|7�߶�:M�����"���0��i�y%�*���nkZ�	j�`��&�i��e�����l� �d�Ϥ"���}�s�8!~n���Mv J��z����
A���ԝ%�K�G/��+�)�|�ЋB�5�"��Ě�'!��)0/�]���\G�
�����w0�ܖ|��L ��V|8N��b���͸Q23� �+X�4�!G6�`ϛ9��) ��H��T=P
x l���Cq�;��@3#�����1J=s�R�T�%7�`+�{�O������R�U? �����]JU��P�&hVp�*;�����Pڙ��eM���0�
8�K�q[���i��k51h�e�|���%L3��Xà���D*���>�c�f�"���FT�0�P��F���4��d�`�w���Y��ם	Z��Ԣ��z/3a�Y�Yy�ƾ[��X������R���P��z�P�PT�fk9���)��Z2����;	o�}4����)s�p��kD����:����Ukp�m��f����I���͋5�M���k+'D�F6=#���K����2�� ������ɵj&�)<-ۭ���?JG���1WZL�-�
R2|��$~\�%ge����	B�D�0���#0����	E�	6�����R�����������m���o��(�>Q9V�
L�>I���,����3E��o�#:��L��J��S0�V|��O�7ɻ�����ŷ���N��'����d�8�6MD�����鲇�1E7�W�Z��@%h�Hޗ�x�RͲ�Ω�`�^Ϫ^��x>��Jmg�r\P:vs2A�A>�M��d��NN��k)#��f�3	Q�"V�ЀT֦גϞa��^�c0�ד�(H�R$h���Ò�4W^���5?]j�撗XK����R�cY�`y���;��'�݉l���`֯�0��ƀ�ߪ{-ؾ.�wTq�DM{��'=����1�n�/�)S������}')s�r���3��ԓ�2d�S���������\W������B��*���%!��RY��kbS2��JF�u-3I��͈z]衍o�a"����;~hH������\����QgV9�y���� ��Ts'����~ˇ���'d� S$�:6@Pe���=�����P�G<�����5�/��0zk����iϪ���e��y�&�S��������LC��KC������JNГ�q|B�%/��y�3��� :�%��"8}��stu[A��~LFX{��UY��o��S�H��5a�pc��W��TC-=8��/���b �08�jL��HrW�܉&q���j2��󵏈��$Ҙ��
\6�������j���#�jIBƉ�^�
 ���ozy�d�R�r�(���)×��u�����O<b�0Y)�la(�f~�����?��D���Զ�B�ն�q���$�����4"���L������70{���,����V,S�H�'�y��-t�gc�Y�=�Ԃ.���{�Cc��_]��3��L��Ԝs$vс�Pe�
�>y��&t�X6p^�-B�a��!�3�0~9a�.�cb�J���L\�[�o�~���S�g���PAw,�̩j��0Γ����%fV�mɶ���!�DC�����pr�7�g	c����t��jؒ�\0���"t�v��	��/-S��y�($F�gU��Vb:03�bat,���<��s�JLԟ@��UC%��9�iK��F�4����f��u�z{��̿�F��Nb��ՙ��jd�)d��eďƿ޾+5��ŨU�:t/F�a.<1nЧ~�� /χ�s����#�58���(�h��cNգ��@EDh��[O���1HMc�.�M>a9|�p��
��j?'����0���vr �Q?���>����n�u}�	�����)˦:���+�տm-GB��ѥc�@�6���XM��zJ�ފi�����l@��1�_���"��^~>5��a�}倎l���m���G�M>�j�R1��(O`Τ���iÀ���p���X�k3e��3�S�����h�oFpYE6����E�bU�V�{��Ԇ��9�Ug��IZx��	&�aE!�<>������3c�Q���|X$���iI+��~���kc�x�z<H��G\�:����nM3�l5��k��W�*�?�9�uM�v�?Sۥ���������ѲZA�"���A /%�`"sv�����`A�B�xT2���|�O����@�����R,�#�;|$��>?��f4��-������S�ڙW�� �5�R�!w`p������q��1�"ٞ��%El���i��Yb���$��k��`$������A{��� ��I�oK�K8
�]�sfZ\W���]��8LX@o��K�t٫���6v<���c2iu�4d�_]��ÕQ�gu��E�r� R�l��y��)$�^e��$�d�� �oN�*�����,Eqn�����HKB�^vԢ.� �����Y����H����T��۳f��C�E�̆_ĄF�|�BSư"@d=_�L}�\(��?W���O)�)�~�L ���2rWYuJ(R>���,�:rH/qڄ��rW�06f�����$����{{�T� ��s��ތ�W���'��,�bw��\*�xЂ[eD�B�2�\ay6I����"�6����J��sh�%]L)?$���}�0�ʦ��>��p�MR��מr۶͜tf[����C|e�}���/�ޭP�CAO_,����B�	/�k2C�~��:�I�����s���"=xww¦����~w�~+�P�m��ۡ�{��90�U��i��{@�#��������a㽅����]��[�����J�)���yčSg���#A��S��'�YT�Hp䵳\�9�mg+(�����R�,d�h=A����E�@/���ԕ)��b���u�T�b_��h+��x�jM�V��T)����e��O�����9�QV&��F�^��w>���y�t�����M���v$%�q�x;����۾�sp'5�!Ը]��� g-bI����2D]a�{%��!�q�&�BF@���SEs�����Ы?��T�?a���G�t�Qf�چF`��6��v�e�6	��1m��K�%���Z�p��I4�?�2�k�j_Z��!{��0��4�0ȝ7�&��\F_[/�$P����F���={}�^�Ƀ̼ �|c����H\D$��5��/\�x��#�4e��D���ud����n&���v($Ϥ���ĩ��~�h�`�?�ȁ5��:>h�+��i ��Q9����a��V�N *�{֔�����Z��l�&Fت+-2='�i�_�B���i�1��R]fS4�dr^����:aA�&R��-����Ƙ�A%2�j�=�N�.��X(���L$��cF�(��  �wW� T0w�\�@G:�h��x�F�H�O�~�������������)@7�Fݐx���!�i��<��.�p��ŝ�>z�j��@�N�����awu~
�9����J��X��r�+�k���D�����^rQ3&s<l��OhhF�a�ruv,)�w�6���E��e��ϫ1)8��d�J� �[�O�`�� u];j{۩�|��D{���'�p���#�?no�����
��df���fa@aQEĜ��ފ��u7���B����ؗ˲2;˿�`ү��#!����^m5�=5�+���V"���w���kV uZ2_B��ܙ� �Pzn��"�K��҃UIi }��1�HJAǋꈅ�D	�/9e�y��Ȅ0ȉU"�N�����9�?e�ˍ�����Q�����@�HT}��^���fIx���(�YH����
��J���lcN��Zz|VJa�j�=�+�d~q�+��4�Z�iН�Fóϸ��>�����9�f�ٓ�)n�P��	R����,ڤ�Z�to�{�!_�&�a?J���U�*�����vݝ�p 5�m)�yIMj~������L���sO�섕y�p��"��ڎ�%����i��>�=Uh2��f��̦/:��I�@�v<�5O��`� ����f&c�����l�;0b�J:�Vt�fl�=�H�����gw`E�"�4��/"�[¦V�(���B��~>M*�]��d���R�r�g�H^G��^�,��~n�Tn�D�}wO{(�0�:��㑄��a軔$�5�o9?t�?D������T8�o���*�$���hB˖��(0;>Ł�@��2����18D��)���]仕�S{R^`/���{��ݥM�ңÖ�VmW���fչ�O�!e*�1P��S��;F�ȶ?���aS~�^j�#�_��L&>3TV���$�"������Q��0��Zt��c��~���q)�!���1
��C=���{��̽^�(H��
a�<�q�;�= tzwj�L�6���{��6��ݿ����F4�<�4(�f�����[�㊹̿.�'���%X ��.N�یr���1T�<p&i����cR~w��gC��Ak2ߕ&�/�cͱ��ye�9�8�'��C�Re�9xAK��惽��-�9X���BsV&3�]}�P1�3^٘��'�5�
��R�7���?_לqq
P�ڧ�>ʇe�HK��O�E��['��/��~����L2��~|5k�x����zefxU#,�3�fu_�H�`�7箚a��ϧa����Av��3���D6 \��J�y��̇�$������p%\�����O �W�K{��Y���9�Q�����&��X
�z�%)�;�<m��N"Q��N{�x��VE27O8�LQ���1����)�`�yz��=�8IV�hƔ�`i��js���5�$$>LW���T1��u��_�X��F!Y���&j;e��H�M6�4��4�w���ī
���Ĺ#"�ċ�`�Mg��oZ�`68Q�����*�#�������m���,��L.3�tE*�l�@�)u9.�4�Ƣ���5�o^q��_���C������(3�'�	�ȅ��#+ۢ�Үػ���F��	9	
|N?���~��Y����¬|���*D俦Յ��gy2ą���gA"@Qmy/�ÝNh���$0��Zg��:�a��b��������,zT��\h@<�m�x2�cRkFk-h�G��n�vᄢ�M�V~��0?���,��AP����v,Q���FW��'}ա����`�$d;�I�a�>t؉�֥�^� @w��w�C%���V�+�ݟ��Q�q�����M�E��`�Ί`�,�{�Y}��M����[��0����(N��H,H��|����c䏿m*�I=�pB���,-K ���?L+q�ƣ�E���!��γ�5�Y��$���v_�Ĵ�������)?��/��+�����*�����Z=��d��0����/I�&i2Ž{�r%OC^D?��m
�6��n��g*ojh�Ѵ��b�Z�$o�$x? �H)�1]i���Td�+1����R����]�c��=bT��؛�ttu��R�}�b����^��=gO�b��*]���Yp�g��ş㤗1�t�!����K���BZ�ݑ��<7��mz#��,E�R%7�2��[</S�)��$U��E��=�����\pģ�0q���-����$�x(�z��>�#E�֌�/*�f�Գ�A}<���|'>���;����j��N��<�!r�'��Iw�e͵-�$Id|фB��� ���fX8�@���[�0,�[[�vB�BQ��Ul��u&�o�Gů!9f��;;-Z�Ҩ��ǣҿ��Ī��r� L���3�a�-���o�-�}}J�`<b��1#s"���9	yi� S����	]�d�^>�%d�?�n �/%�j���&���c'�-�,8�p_Є�����+�F�� ���kI=fy����`Y�d��U$`�)�>�/@�y���J�U����:ʓLy�@����rK5b F/�_�_U��J�%���[��.ڕu3�����D 1�koX��}�-w,6.�����z���?Ĭ}R$���bZ���4������P��2��.����� ����C�97��<�1nߣ���6�~���"�^�,����"3,�@���'ˠA�����x��I!υ��] �Y;��)� ǽ���4$����Cu���5h(�����M���S�SǠ�iJ7���^ag�D��MU9b�w{��P�#�oS�0�2UC���Q�{�Hi��%��Z��$�lO��xa>�F�y[���3���b��b;B.���hw����|�8!i��(1,�3��̬h�����O�m��c#2Ǎ�ƾ~%êº@:��h����U�͸�Nk�{bp�|��g��:�ge�݊��p�O�_�^�u$S��@#H��Y~[7Gx/�ݪoU��B�$B��"�6��\qi�DX$U�G�F�U��c`C���5֔c��8�`�����L1aʙ�?����y6���$� *2��7N.��څ���"F<*Ǌ�W�f��m��'��N���>����b���S�@(m���@E�i�fa�^�w�]��V�-�L�a��P��Ѓ-r������Ez��F+�T�8<��A��+�k�	iw�+lI�Hf$�h�'C+ӌM7.�%�	�(�B��ɭ�fP3@�K�e%�^��PK9m(M+[�7�-4�@�+�Gd�&)��5�a\F{,%
����95��qB�l-ifP��!�o��o�{t���Ѽ�A(s�#�x>1�C�����?��� ��
�X{�>_K�ܼ�ѰuE����	W�4��7]=ü���%`�C5j�A��5�Ef1 D��'�1Dc���ffL��-4G�N�+���}Vk���U��_[��S�)��{>�\����Lw	�Gc�c{3F3Ϙ����!/�&@��s8ƻ�s4��Zc��f��/��%����zs���RL����N�F�7�ѻ��\�Ju���������m1�4���m����HysY:���|%Y n	W&��%.���3e�D�=|�������B�r)�/!�R�gb�`<�T!H[c�σ��� ��>1���"}��Q�;r�� 0��Z�+Rid�OL�9���+L0Y�[ts�'
x���H��M�1�.?�ǭ�Bg���·��DZ����%�t��{�h���������ɵ�+��iJEN$彚R[5O�uo,���H B�ܤ����s�����e����9Q�0����<�¨�6�fv�ދU�s��C�?1� j$��k��.��u�e©�d-:�:�L-���R�a�I���թ����}MM��F�Kxw�r�+\(�p��W2x����5}��g��3�7}?�5�ʋ4V(��K%͐��w<��|+��V瘗�!���/��;P`!]�'zh��Z��L�-WcXq��ǔŇ�sa&�ҦUGᣣHww�!(T0]d�)�,,��V��B�Zb>]��xa�Q��R�h�9o�W=��z\fj���Z�/w��jl��6Flƌk����-I�X6�e��c�8�u�ZG@�\r�Qw���ֻ��U�;%r����6�fؘL�ŭ���U��yx��*)�����Xf�ț��U�vV�%:�B֔
s9��ȿ~�>W����x��4!a��K�OT@�%ԡo�`f�i�C�����/�iU������q�����W髥^W~��k����qC�<�����۩+58������ы��x7âpԍ+��.�1��~�(�ؕ��NU~���vv������e,��	���	d1�Bi��!��F�����TN�@P�Nү
����o�<{s׆��~��Nc�Qh�Pˊ���B���,^I�,����}��b����u�dώJ-�$U3]�k�~2x�r?��[*��w�.w�M~v�Q�L�@&V�%n�_�*G�����y��ڮ�����	�*ܞ�-Zd3��g�#u��<Zs�j��"�4h�6ǩ#��I��mnֲ�w�0a3Y�|66^��wx*���v%j&w�;;1���2/�[қDl�2te���*>��b��c��uF0@�����uF��#��pR~ޝ��r_�k���΍���.�(���n觙�L�������i�Զ?�SM�%�
ٽ۵�g�
�
����gBʊ�s�Dᅱ�-��S���t�#uU���I��F�������@�|v����/5r% ��xM+�J�ѵ������@cs�u�U7���c=5�������=X�AJ�* p@�lX��x��� �Y�#.r���Q�nl��2�����B�R��!����	����@M���|��堝�t�5y�(�0W�%;�&C�+D��#��fb�(,F%��@K��&ciEZȪv�I~_
C>Ub�.cw��j���|��M�����2��X�d�6f�����6/�~x9g����h���� m��� �7�Cܓ�s���ɟ\��a�L�e�1Y�_5\O��Z����o��XQ�D�u���6�3��i&w�R�[}�؍�{�ന�LpL��T�Iŏ����6� ���|�r���wVABv�-1�Q�c٦ɹ��=���g������#^��:c�i���v�@R%��Eꆩnkq�����x]H�/+Ϡ]ɔc�g����S���M�9ꮿub�Th�^�@���^�$�����R;�z��/�Y���~N�2Q�R	�aF^�N�zKy��J���x�?+���]Ŷ��\��K�^j0)R��R3���%�%���.�Yo��TZi��Ԉ��~��gzդEZ�( ���.9<�N�n5�n�b+�c�Ѣy���L�0�� ���=�3�U�^��C�ymy�������W�M�؇�=����ω��IA��Ǆ#�x�ܥ�\�0��6��2�ӓW7��}����奏�1`�wȶ�������>��7r�I�T�m#?
�%�t2��O?���H��W\Z�o�ڎ]�1�6�l �l��젖��0�)<��`N���Q61?���ݐ�j���0 ��9�Y@z�K�:�ڦ?�o�@)�b�	��
Br��NV�B�A7���v�
�<�m�$E]�̖)�:�`��4��1���u���:}Q�4N��� І�9�I��yؗ=.n\��8E��Y"W%wr�z0�C�Q��z��M�0����O	<�.Z��}q�A�A=�s, �/I]���i�8J��,������MB�1�k�h��cv�(9"(M�U�d�ܠ:�%�Sv����wf6 ��6\~�jj!�����E`���$H�m����=Y$AW�'_ޥH[2�.2%�8Գ@?���x�`����ES�9�+~�-uW��G��R�PH��'�w�`H����ɬ�WVS01�c7�귚^ت���*�@A3 ,�ז�t�YFo���e�c�gY��DzX-�!X
�!�Y�49{��d[V�� �v��+9�6�J��M�����>�0�N`�~<�x�L�]��j�%
Xu(s��R�|]�x{�? ��0�K���B�xg��l��D2H-����q��9C��}!I�$yd&�(^��NDk�z�����2�L$:���;���@W�pQ�0��,[/�"����f�I���#Ǫ{