��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:�Q�z�n2�H�U��θ$ÊaU��mZ�^	��H�5y{.	Y��ͦ[.~H	k��A9����[G���'7!6�ܮ]�o(�T_##Y)��Z���&a�m��-�(�|��Y<�`�|���R�좘D�f*�cYኆ�ͧn6�L���{�-ZH�i����qEe��:r�ŕ��yd�42U�ϼ)L���<0
0�u��*b�?]�O���~Ԛ���h��t�������?�
˞�6Wrv^7!�s�Dn��p��Ig)s�N���������u$�"%�2��-�ĥ�I��0��A�@5K��v�w�C�^[[5;�e]���
_��&�� V<�����C���Ս,2*��\f)�c�ƭ����Y�k�2h�F�#�m�6g�Љ���/7s�STxU4sxF��p�^�͠�?s>�P-XWE͟4�����Y��!A�:R*��)w	�a���TF���z�MҚn�iX|�z8f�P*�鳓3�̷P�'V�$=�(�M�${v�|c��l&��vblፐ䉮�-C=9���g�O��vtl�!�Fu5�a_�u,�
}�����U�\	�5���ś�cu�eb��rҽ?Z�����e��:��w���lT�L��[H/XpO�r`�h޾��
%ث���k�B�8���|��q��;��o-�9V�4<JB��.D��o;?Z*�y�;��
O���r��t��!ь�PK��f���y�K�,a�f�A) �w
H�wT �į9:R2���A��:�׵�h���_�,��Mu�&�}GEf�@aK �<Ľ�Q�;2���	{4�L��jC��yN0s��y��.��:^�W\I��$?�mhS9C'��\9Ӹ*h�fI�{�m�w}����'�M�^!��~��F'��<�>�Q<f1;�@J�l�Hep��(�$4��m3$���X
���	�h�"�,�]�r��\��8�/I�ʺ�Z�U6������` 퉕=�A�H��q�r$�8�%|PA�/yn�&-�ZF�]�~�f�J�r�������(�����Ic������n��C�f�v�c���=��������/߂�x+C0�ʢ�7e�2������V��/��'@����̹�����/�jiG<��_qI�s������ꚼ��Y�Дn��W��Re��ğ}F���o{��tV:T?ibC���r���'p�yT��s�ϔ����ha�an���Wc�[rG��nG��BC��tE�׼�"q��;/��]_�,����X���W[dlÔk���+_����;hRQ��"[��&��tOw' 9?]��3^F�f�j����<�&�OQʴ4�4��0v��ʹ���ΛҞ�F���H�
�c'_	܈�����l��N��n��K�F�G�]��/���Ǌ�.�˶�/L�̍�t�b@l�{�]��{�@'�a|P�����h�DJ`����,B��,	�:|�W��SPJ�6��2 �Ը 	������H^(��`�f��in���.�,^�1�Y������[mA%E(</�,��w�j;�޹�poGL���8!3��-�s�X���7ta�ͧz:���_b�(L	�U��32^�C ��a�q�3� �3�ޅ_��H��ǖ�ImxdEN�0ȚQ�/5ppQ���^w�A{�[�vs�����r6�Y�X�(�����6h���6h��E(�m'nF&��+t��}m�>Y�Lx�[k~J����3i��ߓ�-�z�r�Vq<�`k�I���ߛ}0��z%2^�t�x��.ͪ���2e��Q�Jf.�b�Rn��6�,�X��`�~��hanŶ~���	�a�E�,�s}.K^���'W���w��{�V���� �Wm����j�CD�@�5s"��LR":]�S �;5�_��`zp[��M���
�YH2���l��qM��g��)���Q(8KFVnq�䨱�"�]�H2�Ο;&����P'��C4���D[��`�dW�f�L4��Kg1F�՞_# ��s�Wy-�RE=�~U^�F�#�b�؞)&C� �̉�[����O�wԏA��
�e��Ʊ�\� �Eq����6ѝ��BM���.�8>wK�����:2|N��8Ϡk��p�-���xtE�.��)�W����l�h��x��K��Љ���b&Ց������]��gf�`�/��%Bݞ�,412�)����^Z�lu��6�|`�2�Q�}]�wT�*���� ��Y�=���D'��̖�+ O�����]�g&1R�F�I��/p�2�@�0���Y�1���R�
�p�=�?�f�U@v��9�z'�K�wx�-��G��L�`����̔V��VfqC�Ƈ��դ{�I}�N�;�1$[:�pS�"$���2E	1M$=��c�F�V��e��AP��9ùS�)�)���gI��$3_�Ţ�q(��Bˤ�JfT�r�v���7C�Wj�{�PFf���ޅ�c�����i�����WN�㡖�p�ai�����)��[�f0����co5j�6=��'	�1=���FD�U��<R��W|�l(�
?[��ƀ����5oE�B�<F�~0��Qg9�HN�l���g�F�� lPOj�G���5�����ΩU��7�����.6[�Gq�$Td�G�%��Zz����h�5t�64��>���uA�5�Pht�Yv9h���`}�&��'�A-��'To@�s�-�o"޳7F���ڡi�R�^5���9�V����$�d�4��Mݤ�#�6|�Fw4�Zm�(��;���P�^ ӻ���%��`���xr(��7g�֢�mR�C�4Z��r�8\����8(��wQ����3D7#)
c4���5K4�%SH*�({�cb8��x!�`�`�Dzq��ΓUK�������R�L��ېGw�߉6+f����D8@o%�/�Z%l�R��G@&�$�)Q��
���n(��L�P�7���ND�!�?op #���ʋһ�Z�t�X�βr$D��Ȱ�>J��`��W$%s���ʏ�=yʖ��[��"qcU��>D�Ǯ  H�F���6�t���J��\��9��ń��J�#ѯ5Dxѿh��0�̸B4=�lc�N�}��s�?Np0co�����m���a��8ƴDS�W�-_��ak�z��Aj#Z�5M�L�o��t��,����<zE���I�ի��hE"�Z�wk�qh�`8��#��܎�q�B��$�'hӅ�z���0�ʺ	dJ�\B���r�6j/܆V�ۺӆR�	��s�>8�ќ/�0�,�������Qz-��Y�+�:��k�,˲�.�0W,R���;�cR+�朏���%�U��c`s��`Rj���!,�{\C�꿦C+�Pib�)�P4�M���c�[�z�����@<��TIT�	��kƅ�M����b�:J�m=������"��05��"�h��S@��8'�c�,�L*K��6+V!�T��?}��`�8\���R���0��-�*�8x���?PT������5�s������Tт����D9���|1�$�)�%��'�1\\w|N��p������-E�� j��4����uW#��μY��DU�_��Zk�h��բm�<� hu�(�X9���x�S��[�J�fq�cdȸV�Hi��0��l2����4�30	p��M��O`�F�`3>�U�xJ�B̰gΐm�y��i`���������{N$�W�)k��ژ��K��x�:��-iA�50�N!�;80��ڇ��p�jA7(;6�N���%b�����:Ն3������ܮ!�������O,\�����0�k�����d����N� ��]�e��AJ���L��;�KC[Q	&' �6��B��m|�U�4�8�V-*��|#��#PXJ�%L��חbm����/��~��O{g0���߀����%�N����b�~�徆�4�����`)���~bBW����=�����t�Z�(�]�z*HK"��t�~�V���z��C>&��R������s��1�K�і�W��4ӥ�DN<GX�b-6	�зeG269�+�\]Hu�}�������~��
�8|��� ��0��.��1d�8O8W
Q�c��
�a�ƽ�T-7���M8�CD��!�_8����+����u��&�8 ��9���Ez=-�n�ڣ
��_��i ���]O8R��'I�DANH'|z�Y��ń;h��,�0��3,�ȯȤ��J���*'��B���PF�2G�"��b,��8O�}r�!��0댙�jd�O��ژ�>B�z�9_�SL0ltY��a������i`���G���Ţg:�� ����`�<
v����JE�	��ah�ӫ�2�H��J��G�_[������ϑ6&6��ͺJڮhRc@�gWUy;��z(:L<ˢ�g�d>�������G���\|�fd~��V"h�	�`�Aw�d078��T�N`-�zr$��� d*�Ό�R�!<���]@;�bs1����8�YVL�J�D��M�1�{�\��}�	U]��)�Y~�eSu�k"����Y&^���{j���M����<X���20]g���5	6Z�tFm���	}�����g�L�&TI�/��g�2/�v5e
�&'��+v9��hg��9��σU"z	��j������ʕ6�[�YA7:تe�@���J`ZifK����iOFx(��Z���Kv�Bo�C���t�<�Ͱ��)c~y�r�A�x���P���mDn{簶��]�V�����/��:_���R�*����b���GGVcXV�.iu��\z{��4�1�F������Z�GF��i]�P�=�'��@S�!�Or�u(.:#��f��-ٻ^���Q�Љ�7,W��}�ĕ�cX�Ǎ��BR���z�8}�Ĝ����0}�sDJ��a�[������ Qc��J��/��	�Zʔrۏ��L��w���W���qi!9<B�����"�!�/p�kv-��XD%�����k����US����	�>F:xI�$W���tA-�����&�y�8o�S�)�WN}�q-����q`� ��j+�dk4��K�/625Cid�X�WT�\-��D`1.b{䔪o�� r�e��ܝ��.&c��qh���}X29O@���7�Z�����Y�����>E�|^*7��a���e�4�R��*�`�Ǻ�Zc��,�@(ˍ�s�*%1�[�.~úi�Sw�10����uG�݆�*���{@��r��`��~⚛X=��¡%�������T���h[J�T��C
U���In��õÔ��l����]�x1�"xE�G���#�vY�����[h!����?�E� u��|��.�9'�V
��v���0G {��&d2��=���sA���@fҜ����d�XR�d�z�U#<�G��i#d��}�LC�P�r��~�c���|UG�ׯ?ig=�r�|�x�W��|Xx�o�|hsJ��u`��bk^�j&�w�f�`�װV���ː�sm�Մ��ӟ��f�a�����������讌�����Թ�ˍ
�5�!|�g/3T�i9,]��{gƃ*+	X�?(����n��یhD��r䊂�]Lo��yr<≫c[-t��,�S���C}K-�q��4�7x�!MӺ3�wW h���-�NW��)OtY���Tc:�j�DsU�����$��l����<����1���Ҳɥ���86v)<�Է�G6�_3SS�F�t�������a W���R��N�n3*�=y�MS]�F��!��ˀ���;�n�Mw�u���U���Z���U��Z;?c���9�'���U4,���%u���i �_��WrEd�������nԮ�=�m�я3�	��y�z��d��)<����ѫ���7�ԣ��|�+�� m�@y�!o#�@6��:��U��DҺ��eŹ}&�\pH'U�N�67�3�o�N�S*6���&�l��F����i1�dw8W�q0�`p�рf2�	he�p�.�E^�'-�W���qO$���i*&o9L�ˑlC�7�߯R�̙�L�(�=f8�F:��D�;�t	몦H�����7]Y�)����{���箊Ix΂��<ߙ�٢�ۧ�o0�KC�EP�=���M�eiY~��80���̤S�|m/�>�X?���l_V8������<|�]��u��hO��9ܜ6����? 1�a(aX8E��44R�����[5Ċ�o?D� ��ˊ�m�������~n�{"I~�TT�z˺p)�.���%]�*e�!m;�]�oP��/�h]X��>!�{�����&>�����Y�o^ڽ���a������c�N�5�Jq��SoThK�ϣ:�J�]0L�_�Z5�Z���x�mrh)0���Do�yga�Η�*�6.T��d�l���U�/���vq��`�X�T��aߵ���>�W�$���2D^�-���YTv�L$���\�߂'>y��VE3��5J\�Ƚ9��D�/!3�Rm���_ʱ�Q!�^��o�!렔�6�6�,8��n�t�ݮ9s����:��l"�Xwf�F�q��V�R���>ho뿳muDB���\@��tr�����fby;ee�B_��uB��y����W{@̛$L"�+��[�\go��i��!�F;�%�S���+H�i~�M�#�\�!�����?t6Q1�U]���@T�%�0&+�^E����Xn���z�}�on]��SV()k�I�s:�{�.���R�)��YQ<g��D�,N�V�m��υ]AN_�|˹uҦ���]$^y�l`��@X	�r�_����a�]�{�iB�fm;
ʛ���U3��K��N�@�`M�|.�k]z�Dיt��U&v�u�D��@	���-��������DcR!ئ�#�Ē�}3��6�A��+�W��5$��~�Ηdx��`@��-�|=�~y���k
X���W��r���]��)/��@(�&��幃X��p'����r�n���7��5�ߪ�J�D�"2�"p6x0�fV��Dq{�n���}�;�}֬�h�����!V��]��ΦH�T�R�����OEA��F�8�5�~_��@§�XW��\a��b܍������]⿖	9=��^�}P ) ��Ɨ[g�_-GQ-�6߾jGQ;s�#<��r�Z�$���`�/`\0�(�ܸ�'iU���.�$�<�#uks�����b��&
1�^�}��u��5�x��.�Ao�'�˂O,��扳I.v?��=��=���$*I,�O�.�>�hQ]��������|"��2Y�����I1�4dFr\9��U�<��u%Q;��U��Z�S�4��x��W����g�7��g���X
�KN��k"��O��E-�~����md��D��w��H뇮�g�5�:<�4p�u���n�װ��m���.[�a@|��\�nQ)T;��
h	/�����<�$�]�|)�RU(��b�x3�Ô�o���ׂ@k� �M����1I�a�-Evg�;�4jm�0��j���?��?�<�G_Nt�j����t�.��'�/�c�#��� /�!�ɒ�NCz�U5�<�[ە�A�߂�^��c�^�8-#4�Ha��~\4�|��E��t;�q�m'[����KdFzn���ى3ۯǄ�M[��{#4��c����o�:��ţ"SY���{�$-u`�fƉ�1;���@j�?�G<�K�zE&��͢�}��/���/X��4t����Ӌ�ּܐ�a�=�H`�/+��зU[-G��	�nf#���Q���3�✍ �<�,�wpvK
Yʾc/�����Gf�A����QSiT�*k:���B�dw�]�<���p�?F	�~�:��ą!�މ��9F��C7%�ɰH'c,�,�9��/���k:���	A_
��]r�:�hmԾj�d���y\��:��ps9p'�1��0R�*)��2q��K����d"�=0������Q��g���2��҉ h���Bf�2o��ͅ��m%�3�7��{�Y�E g�G�
An^pS��J��p�flL��|E#J�{��p[����+psVA�v�}��q����6Б=�7��~(��L�˩s�Ee���C5G�cr]��S�/��9��/J�_l7#~���;���O!3���p��:;G��6h�OAL�o���ιX�l1�nX懜KUB��*�x@�b��*�(�����KlDa��`�n+@���X�+��f��T���,�5�<�q�_٨�V`x�Q,�p8w�kʺ�m��&�k���E�Y��q���n66.�j��؅�� "絾�mi��"��8V���׊��P�\���&��˰] K�+�}��u�u�f������(���[��'l�:��ik=��c����nR���&j8c�
�Jd�Z�������ê���r/�+���]��r
��$�gϠ���Ѷ��ޡ���ft�G�m���/�(ґ�Z�7�=0>'��R��j�D���m�j����r2���r���פ��JZ`Idc?+?#	)�pM��E<�td[�@~4]+X�ʋ)χ���g&�*�ư���c$�k�I���@���Y]ר�g�."m�U�3(�Rs�0�%��I<'	�S�K�I��˅�
�룛댓
F���g�p�Y���S�/.&ҽ�\-� ���|�gz�\�$[��GDm|�|�1�-��`U���(�8��A�E������v���ƝѲ��ʷ<�����Y��YOj��qU�5 ��sO�ģ��w�w�~|D��^���.��ˁ+��H�n�L��/'v$~����ݗo��V�ƌ�����ј����i�V�*�iv½�AT�8�����,����{���)gOG3v�����5�n��"Rˑ���B"���>/����R��_��θ�AR%���w]Ԃ��9J\���,ڊ;Mq�#P�q٪A��8��$�/�p��d[pT�=�J�~��9<S�9�t�y���RVzȮ����<�bh��F�#ѹ����	����R`kx���o�H�����m@�������O�-ۢ�o0�	�WL#V�x�߻j��5|A�[ln����zEEϦ����kq����������������%�1Z��KO�G. ���2���o���D�Y���Nْ������f�a0�=�ȍ#�)^�Ur��]� }.�|K/r� ��^������@���Mq��3���,
d�_���>o�+�Cz��Qs&)��U�%խ�늫��Y��1ݓ���rc�#��еA�
\вT�h�Z��":��<5(_V�-ʑ[mBWJ�U�}��m�P:k�o���q0/�9�R8~q9{k�fCΘt!���ug?�e!I�ڻ��|�%f�}rT�j�Fp�|wα T��Lv���s��1��WeVR�`p�(cP9��\oK��gʪ������h���#��H�5�a�'Z�v���{���R,�f���I=���M|mO؀��tT���F�>le0�Yh6a�X��2cD��/�*'�֫��'nśk?�]Do�H؜�%�*�|:���
I|���\M (����s����%o�hѠ
��ڻ��>=f�v�%ۙ��J�/�\�3�. ��[��Vu��(�ײ6Tz:�����2�*���i�Z��D&m[P�"���_50�kPz݊6�<�[�hT��Ԥ$��G�C�&�ڏ�_��SjZ��v�\_���E�P^�eg��ʬs��7�f�]|��8���і�΢��;��F�{�������c@�D��r ��ݢ��39^W��@��cM}Ä��Q:%x�^�j�k-]��Ũ��o�w�r�7ռ�40�*_���I�R�Q	k��HL�tL������
ܒ��lA*����W(x�1��~�RN�_�np�AQ�8��8����zϿ���*���2���޹^VP�n�䛙�c�rɸ?��kj�"H�} �l0&�*��.��tY>�"�<`��m� �=D�%�@J������R�";K�B��s���cH������� ��\,��?��6x�v�V0kxT?�7���H���T�����vN�p�����r�Z~�z�A2~4���t�O�
�J�<H{�nt��ߓ���&�u�'�
����|@$P��-��5�i�ZwL±�����:�����x�v!1xW�)8�s@⏦" p]j5������B,v�݇���{x*Zb	�M��*�<B�B]f��w�F>�\MG|p��n��͆v��b�Z��K=�{ǫ#�����&��&���ɾ���>tmA.֨ ��Y�f������I�Þ������Z�w�'���ʜ?U���,��Zn�-1"�S��D����%�/���E�K�8��:&��҄�(�@b"���?Z�M_�H��̌o+���Vz��y<��`�@o%�5^�-+��(�M��k/�;���?'ށ��p�����V5GVM���`5���eyP�����;@�$��%��k!�!P�.��w��``��a��[��gJb��G����&VDY���U1��	�Β�%d������Jx����/g+���p�;�̾pSO�1���j���sq�b��*�?R<3k!������C��������]�Pj;w�v!KRE��������)L�2��*�����E�W�jkP?z�;�ԯ/�H�s�ZJ�o懗#��U�f9�3-jǑ7:l@�:|�f��IYJؿ�Lݝ��X��l�k|����c
���<�l�[�u �-!�\w�,٘���������[Ȑ��l����(��;X��~�O��(�פȞ��~rIo� ���Fe�)�oZ3��S�>�!�4]�h'�׻s�e͜"c�����{;�!�g�����Q_��L4yI�
,q���%�:�#����Hx�M�&�E/�Ia���q1��	����Z-d�� 3�P��&�mj�%�ݔ����E1��%R,�f5��7q��n�aƹk4e�'���y�$d�<5��V��e��w��B��qX��T���d
wcw�h�~(�3�y؊)�	&����
��j�U)ח��&��H�\/��^��>�ef���pO�_�Q	�@�'u+ͱ�E���!����%4����5$:f�
a�x��xg�;�;<f���j���wn^y�[��~G� z������3����-��h�O2�FBT���q�}xD��xO"��9���������c��i:�Vo ��ч5Rj��W��[�O�_>��{����S����oG��
<!�Q�k�G�w( �LH�܆�ðܖІ���e�?�t��Fy��Ս���_��ԡ]ֶ���h��?W�
��p#�N��h�q����ȝ ��:��C��Q���BH��yfH�~�&�6��KðQ�Ɓe�� ���CO�3��+���r��i�2���=;�Gȗ
�!�_�زy����Z�γ�/�?=����ez`��9@<�7� ��XU����u���{�����в���c)�M
��sthG�w�z	G��2���wU�<�x��Bl;ҙ�`%���;1Θ�c�h�L�z�� ��Y��q�uI{�D�I&��.�J#�F���IeJqyfYO��qVU���I �X/ـ��·lp[ly�&��D��F�8���. �e[��Y�K��A��V7ua��C��p����]��허�H���m�A�T��vASQ�DY���쵖�謳$&�@l��ȒJ�أ;%R���珣�/�׃9��]�>P���yjF����ʽd�"�@q�߻c\�QXTЏ��O�{�{zWW{`�>�n'�&�w:�LRͦyp奇8�wo�a�f���a@�yP{\e�d���2�b�%��>�&��z)���N���ϕ�"�2�!��S��G�;D��ݍF�}!��^�ț<e�����TLok�p6s�8��1��)yiZ~����g���}�k%�r�m��m:}9��`�Z<��)K�ZO��+��� ����i"�����̚poR��p|ʝQ�3-'wt`z�υJ�;��?�b��
�EI���)�e+�4P�Q͔��]w@̬�]�ؼ�Ebxt���
9"0cHy�������O3�uP�}� ��v�����-�3U��K��κ�W	r5�Y 3������M�}�|xT�˔'�3@�9�(�D���YL�`�&uo�����4e�!�;	p!��~�a�\�;0A�'����b
�pPd��Y��j�H^?/�sc~�J0�Z{�U
��aP��ό��
>)}fmE�(��*��B��sy��"�xB��$�-&��@���\�uѺ�^򕖕P��6;��F���9� H2 �G��xw|�^&`Xv_��А� ؿ>�8��4��I��\���M���$��d���ڵR�B'Sb�VL�;1�	�+���N�����m�,�ɚ����{V��8�ʳ�K@��&g�G2X��L\�;!�8�a����tK�O��������MB���/��O�Q7�9��� s�5׌���Y�TG�9o�Z��4���Z�
!�Ҹ1���=�@2ҳr����޻��*�7ĩp5�KD��ÕU9�I6�?DN�;H��Oe@�p���K��6�� ��(���	CW�)��}��W7|�J���ޔ�vGT�ѯ �!�b�����0Ӳ���8���]�q	���������yM�S��c�6��h����`6�����҄�v��r�=M���ٶ��]��|�Z���+9Q�>B��ap��2㡤��ur�(r����k_I�\��?ں��BYT�|أ�}���8�:�-�)�K&k�VYS�40�,��t�n�}5R�i9aO�s��1f��Had�o�,S9��;=��A>�2Y7b�-Т�3Y�G�%��<�_�?|�D����x=�R��c&��Hj�巃N�e.Wj��'��] �[�Z5$�h�J����y��|�j�k�C]���{ٳ93 "��hf�9�e�}��S�/��F�GJ�3!DGZ��0�sa�ñ��~6���HQ�t�| ׷��/���`�fmb����ex�?�lAf�e�] ��b6�w���}�D�R�t6t�����j_Y���/FC�
p	��/]#�@�a�JW�^vbX"q��su�����(���=��3z UY����$��wF�q��x�������,"ŕ����h��Vv��T}�`��!K���
��v��	 Em�O�czaׁ	Ed�>q�F��-Ӣ^�����c7�N�dM· m?�-3bR�*K��a,�5�#�=��w7�'�#�	��d����<�$+�&D��G�[�K+FwgVmW^$�\fC��~��bW���6�pNR�+�:}	`���i�ϲ��y�XX��i�;GD�3IO��H�Xy)��o>�H�G���,����>@��i�6�4��7$�_�.���զ,�qb��U@�.���s�����XA�J+��5�u�p�*�o#�2;��K��f �Y��G��~�6t}�U4���~E"�6$i�g�"w/z�ݮ&Q �G��R����Aן���_� �4V� :C莊Y��ܫ&��J���6|��E���b�(<��nw	MK��c��8�������T�(=@_ʯ1�ɷk���-���4.��B[F�{FE�~I�i�"1j�'�V���T&9qN)f%�>��u�D�۲T�ߔ�V�}l@�ĳ�ܵ����~FG�+�>XU�g?xn(�am-�Q������h�nd�IU�p߀�����<�כY���L���9V/��D�M^�|(��ɉD@E�#��UY¶i{sG�:�xS����~!�Ш�����MC�)mOؗ1�.U�D�H�6֐g�l��l=N��e��|_$�+~W!n,>çbx� ��a$�'4��z�s�i���O�y��~g��s��q�G�d}Qǯ\�wu;7O�tedC+q�aD��~��h���{�:���6������ѩAN��4�����}b~*1��d3^$������؜�9��o�w������]M-�s|�9U��,��x%Cej��E�-��(������xt#����ڊ���h:1��F�}E���m{,ۗ�\5j�����IR��ud��㜕Ӵg\��9	� �c0q�E���`O<�J�_�P?�-.
}�YD)޷�vƃ�0�s:���2��.�C�N��
}lwU�D��^��@m��jòt��lÈВz�b���M�a>RV��3���,~�j1nl'>_u�Z�mM��s�����A�mx�0r��@y����R-�(0��}�-]���g����̰ᆜh{��@�<n⮛��
����T��9cU�<?�	�H�M]x��/�4�7ql�\!�,V9(; �cWI[+vn��:�(>o}Q�^4�������]P���88�5ߗ\�;1�O<8hb��m��Ѡ�a�D��!�۫��Kz�+O(;-˭4�%=T����}s�6��T��>�,��ܳ6� �Yz��]J������v;E�~�� Ϋ\�+���F� �r�)35M@Ԫ�
ƙ��9�P��I����"і��3�2ǅ �Z����D��0.!�3T-vE���Ot�Sk��L��;�`B����m�@�C��!�8��[�8��8���m���P�<��X����C|��<O_��I�Wx��E���k߆#��7���`���9�\��J����[��(g�J����� �|�#-Q�9נ��&�����P��Á�p8ÉIu�_����0�x�^� �a�	�W2�C:O[�����A��3�Z)������Qy��Q�H�;�������b��ͪj6:L>]Q�:�"����̞���-�K�1��5�hA݇�Xʀ"�.��*hu
!�3�c�_f%�����\���SXc���Ƨ#jF��2�B���v�Ug�6sgO�ce5Ir(��a���I��F�(5�^$�X!��
*�(
%K��\�P� ����]�+�9�ɬ��$���� �V����Ѥg0��)@A��E���W5�]]7�׿qZ���ZL
�sV���V��!)���CD�N}���;�v/�4��#����ݿ��\`�m���`�s��,�����U�����P��E�<��P���8�a��ر�6x��I�� �����J�@ANb'.�͏�I��{)�8 ���k�Vn~�`�7���K�HQ����O+gE?]��)����eqc��`y^Z�.��ҙ��Ke���j�����@���K�R�����4�G�ઞ@��ҩ�q[,!�����=S�%�ol|�ʽ�Y8F�ۺd�k�nD`�Cy�s��C�;W�_�U[�m�ͻ��2{������g�T��#��d�eE(w�ꐔ\�F�ྸ!��%t~�;AG� �����$K�����y��T��?���2��Dm��ӛ98���_������4�f����j��װ���£��;��e>Ov6�j�0H����@
C��e`e{��.xh�[vd�0D����+>	������'��Xp@�8m!KUPoˀ��D~�5���_���,��u��|g0������:�ab}o��؜aG�z�Yx�(ҁ���L͎�9���3Q�;�
���vT�sV�X,��s:\(u*N�x��E�ӿ]IN+�l��+o6�bP.&���U]�D�͵��=�2?�L�"�g� ��h=��ښ���as�T�!� L��d��z�ա�tՄ�s���=����lF�
s�s������}л*��0;e]�o]1���!Wo`]�Z�s�GW�<�[*�g�Qΐrt�ӣ,���6�$"��?����<Ж��|�ԭ�	^��js�^�d3��*`���]����p�HJ\���64���Y��~F��t�t��>�n��	��V^����0��o=�;*��;�<������k�+��/Y'�T\¯��t=~��l��q6=G�&z�	���[���t���a曖�B������f_��ݡ�W9�����5�)`��Q�۶l���������>��t�Sd�igE�`i�f�?潍l�r(%<"��[ӷ懲6#�{G��	F��J�Jv���3��r&'I���f�6���k%�4J]�]�e1(�{�m��'B|�xK/��q?Jt|��������g���n�}�9TO�pi�KR��[���ټ&�&�_��8��
gn�}��� ��]N�-[�Z� �o@�fa�KH��ӤK
bi�G3f3�mF�9\���vV5� �$"w.-���|r����ՕR�q�W�S�F1���q�����9 DJ�e��{qKm�X��g(�$��n�R�nج"Z�g�@v�k�I���>�d7�-*q�M��مS�F����:�0><z��I�#��뽛F�AI�[�q���f�	�8��>�̄�W5�Y����v�LE9FR��l�f$��Ia?eC�����eu �.{�C��w��� �
c�ءǺ�tu������8�5:�[2�l��!�ctj�4�*Ic�U��Y����pi[��I[��*Jt��B��@�暇�8v�"3i��o���w��R鿦�\���Or���S<�f��0[h�!j���I>����Ik�Lf
2�w���Ϫt��H8
���g�r��-W>�s�}x+�m٩>�X���*�s)"��l7v���M�k�+��9�s i��ƌG����B��K˴���`�l�Q���ߐ��(zfa �wvl�U
)B��1o*��6�Ą�f�P�ѷ~��)�q?��z+K�SE��G��~%~�2 Z�6�t(���mR���`��A��#��*��eM�fv���.���+�a:��Ҡ�8�����S��̫�ćY����[B�Rήź4ځ��#�k�^t�Rv�9�	���;%��ͽʏǝ���������z2q�첉���u�*Ivn�ët��ܹx���:�FAȃ��*����"��F �R���k�B�G��D,��������R���ּ��Kd2���C�����J,��������B+��L��F|h�i:�9U58m��:N�%�F�}�E#a+�$�a=C����il�mu�c�|�Lҹj��Wi�h�:U�'HuʞlQ-A�$���|#��̿�4*�6��kZ{(���F����쯴���!��A�&�u�*��?`��2X�l��t�iĲ���+��׻��U!(i����"�U�����L��#�%�����tjǯ������f"�-��kT���:��O���0�������;i��/5+�c&��d$-]�9zR)ͥ}�d��>�&��a�2�Y^���nm��>N��� �U������D�J�=�ԅ8�Y$��Ql��N�+��C�#r*�*nxЦ�"ls� ��5�i;9�i��rZ�(s�BJ�8�����-V�P��g3p6϶ϖ_�����[�CՄ�Q1�M�y���qjM(��;���7g Lɾ�3�؃2C�y1袭�8���iM�N{P�2�0�k����~ba�o 3_��:X����o~Ko�4])�k�6��_�;F� M�`9��#e���+q��/����4B暄w˸��\�g0���d���cEh�܏=R_"��Z
KgA��*�L�^3+�|6E^k�k����1}�f���i)�]�Єr��	�-�a��JE��-�rǍ���M�m-��A�f��Y7�pGu����9��D�KRM3H��'
gI\@��[���4.{�&�^�y�o{�����mP��k�$|�)3_4T���Q�D&���@<<̐?���~Aʨ��ŀHu�����۽�Rʀ�p����z��
�9�����D����z�F�SD^�w�B:C���A�s��%ds��X&�ʡ�A���+b=�#�=�G2sU����p#�=�]F/���yM���eדEt�_?���(�.��^;8�e�1�X �/-�xZX&���s�H�����F�b|�)����Tq��p|������Tf��a��[�Fj��:��1E*�PiB������@���q(çs��h8��l����7��q����S|���Q���K����y��Ȉ~�𢆜�U�sz��H%�r��M�1u��ir��R��.Mr�K��Q��ɷMF��>Z0O&T��v���A9�&��S4E)/��ǍD��z��'�`���y [W�%w�7޳A��5	�:���[�M{@�*��R,�-��Ȃ$za[��ʽl$UU���C��K2�x�,���P[��'�M՘u9��:O˹,�!>�I�9�6G���q	ʺ�Ŏ�-4������wp�$��X�<H�@tx+LDe������]���S�c����9w��97�%,�x>��R����@���-����a����Q�0�k��3����=�b�];\8�j�����0�m�k�̦u��摕*x��� ;�]�IF�eP+.�ܬ��Ǻ��J��?���0��d�뒶�+���ż��P����}��k5Q�/^kc�0wv�G�1Q4�n�����K�����c\��S (D`}�1�v��������$�#ё/��������'�=!θ�\���cJ%�*Eq2\�a�V�*� p����Ax�yq/�[]��axif�����NG�c�\^��������k�(�ؼQd0[�¶�:��ŵa��x1?n	o.���C�����O��3t�y1.�f�[`V��o�B ?N�. ��ACv��H�R����A���o�}��P/|�/�$���@|^A�[��p�@��HP
�GJ~��b����l��Tn�Ff�f��-9���\q�	�B� W;r���8��ݪ:|Jk�j!����"�����o�\�>E�H��\��P�[�.����2궗��K���ݲ�q���WJ���=Ɛ���x'�o�	E���?K�a;[9m�(�F���Yp�|�m��@��
�F�Ŗ^#6����Z�0��k20#�h[-�	!z�*�t�\���2��uyq����  ֑YQg8� R٭ߓq��8~*�|E4
pq.T*l�b�zv�!�1%��"{+3U/�
��n��H9�|�ɀ�ÛJvո?U��a$f״M��3QX��;��t)3%�_HR,�X!������p�l����jB��.��a�kvL����5}�->w��ⴊ�P���L9Z�5�$��9���Pp'*���S���-�=��spIRN�E���>����⎭c��p��tZ�����@�(ǘB??"�������N�~D}E�����[�,*�`���YJ'�~���4r&K�6���t�甪1��n���[�Y�yMGe��Z���e?��^g!(���l�A錣`�L���T?)>�\>�.Z�.k�A|�rz���~ ��51 :��"�P2W� _k���ʭ	������i7
X*c���h�����]dd�pA�D'�j��7�9�E�4�Ԝ��O�7��e�؋�~C��i^Ю�½um@�ѐ�5����K������� F�2�5�����*�}y��M?]�9׾�op�ԎȥN��aa�ڞ�3�B���� 0W(�&0�s����/�k����+ժ¹+��e�L����H�$����Q1�Q�,&���-&��ҼN*��(B�Pl�����|qhI*3�e`n)3�v�dl1�`�<;p�B>T��蘿�1����ܮ���q�u��Y�&� �Z5!�ۙ��f]�w�T=z$�{����g�QUMS�=n6�'���D�~�6Z�G��HiK��f��9O���Q��m%���[������-����6L?͎N�s�z)�G\���� 0�aӮ���\�@�B�@��)`�=/ ��*Vz�/�.�>�xb���h�V�TaB?�t�8����dP,�}�B��-���$�Ϧ�̈ʁ�Θ}z��	=Ny��l�KX�����~�h
\Кi�E�6���f Ϩ3on�����rp\A��B*ra(gk�pf���)��P�zR�c���*B��"ǓԼ���{w��m��E�}o+��g�5/(Z�Ŗ����B�ŗ	5'@��T䉨�C�;�d&~3���Y9�D�M�7�IB�$���O9���8Y���k�G�L��Z2}�.�-��T�Q4�2�̍�TAJr:��ȴ.��$y�Dc"��Fef�q��@�u�k�.;EwD�?�X`oP�V*]����HJzfo֕m�p�$��&Aua^�f��Qa�S�X˧ �<婐�:FtGz�B��Ȫ��򄟻G����%$/���H������}���x�����aDRng�# ���Y��e��Q�o�9�o|}�'p4�msd�ƒƱ����3�\4�G�X��%Dl�N!}!���~��6� j(W}���dgx��!C�RZ/�u*���=�Awr�B�t�_���'�ؼ^��4~��oSN|���Ct�/<?��9/\�Fk�#�L���B�����K�y�2�5m�8ː^�]qw���۞K��s{C�d�DΑ��_�ӒW��(�(>e+���h�����S���z���#?�%&�@
�l-*\E5�x�r�L�zqMKxa
�Y���W�S~)���7I�����{��|0,1h�2~A;v��u��HO�0�ҫ\���"(�(�Ĵ�K>��^�|P��mW����1�d�b�=�K)��v.�u%��U+A���Q���I�3>��l�~[Ҿ��9�c����b��;����M=�Y9zl�d`���7=[��TG3�	6DY1k�	ݸ)��2ic� ��3���@Wc��gO+|�&|��p�y�������l(}�J�PZ�z����3�Pe�o��[g����6��|�
�P����2I5� 4���y`na���}
�	��u@��e�qO6�L�1Sw��o���
I��6��[�
W*2�}�_�q�kE5�V��?��/�:�G�>q�����T�7Q���,����Wb,��Pl!�� �3q4$��x+�O�N�c�d3t�Ez�b�G��8���̥Ѻ��mx�h�n,&
q�2�%i�G�:|H���& ��;(P��[<�J���-!J���\@'����z��߇[� �䳬�L��<oef���"n��n��Rp�8:sW,3c��@�����E��DjVg��Og�^H��X8x(9Ʈ]*�� ���b�;�_��ԐA�,����Ns���K��>�?���A`j%���1���(�ϔ��{S]�����@aJ�N��D�j�+�aڏ��Mx+��nR��v��ʑ)fŋ�_�%��	Ѹ�;au�G�7�� �N>R&,vR}FR�~�\l�R+*$��$;ڍ����2�a�r�y����d�d�ň?9������CQ�ɣ�=�W��ب��=ObC)x�#������y���g�@����0fl���70!�<�$>�bE�p1�3	o��(�'����_B`CP��;ݥq��59�*�;�����L��u7}�`LZ �)/x�I�1XU8)U�={�,m�<���ZMʔ�d����G�|�c�L�_��1C��J~��:tJ=�f���O��ـ���&/&�yy��F A�oT�����@\�q㘛L$g�
�DQ�Z$��ªp85A!Y�k4o'����L+4C�VB{n����;�oϠS���
�v��$��D�t������FLW	�5�g�������	���Ԓw���������	��A�}𯾯4e�}������yeZ^+>��V�{Z�~�Ė�P+����t��)+RӚ~{� в�ޢ�= ���t�J��`&Z����}����[|-8Ǎ}�^h�k�GtKC�R�H���\~H���I�pr����^2xy�v�er��׵I�'fU�C���at�^|D6m�ؽ�����Y"E�6�;!���6;cv�?�>� '^�&�,����%�P��S}d��}H��'���Թ����(��{���e
_ĿK�e�"����i��ĉ�Q�#6����c� 4�·�\�372�+���G�*28���CV���`����S��7u�b�ǳb���E�wA���p����C3��SD^๥���6�P ���	s?FT�R�-�;M\e�ؚ����?Ǭ�(۴Y��(�ؔQ���#7MY=�2XMh9�����<f�0���5��|!@��"��ø���z�r���Fc�Ȑ^�+(�������j8"� .�K��S2"�bt�ꜽ��D�=��f�Eh��mk�k�ڭ��$�@�%�J�<.L��G*�i��u�X�nnWW"̞����e1Sf�A|�#�5IE{k�>����
Y�t�l()~���?�rVFV FM�۞C�S�b�Ɓ�DS���A�X�����h����|�ɏc!�i�-녛P[�
���W��rt���S��n|�8�����,��r7i��r����RMχJ=w�"�\��aaK���Gb��b��>����9�zJj�(����q��/�x�<���׏�|���o���F���q^8��6+*r��cf��3����i>��b߆��z�'���_��i4oÜX��2I��U�ΉlBtv~��%Y�(��� ����fq<�}a�Fh(�l�϶$QS�C�g����tT��vS�u��)�8�ޮ��-�����!����=���#
��Uc;�K��;׻�*ɰd�ո^�Yq��Ǥ��U�j�F�|��\�}�1jBT��'&Z���{��E}h�X�f�p�*Z$T��LB����C��C����� �p�6 ��kL���Z6����W����U�,z�iywkl\�c�[�˲&�3l,*��A��:�C2ݐ��7`�s3�4i=����K^��  V_�=4�V\��s?W�^:h�<�&�1�\��.l�nn~h�{6k�̥��t���*/���|5�4�� ��Üv�|�r>����KRɵe0������B���zA`�y���nc��CP�f�$తR�_N�E��7���H�*B$�i
i;�(��J�ׯl��W2F� <�}t�ru�/fVXu��_�[DD��Ţŏm�a V¼��nn�x4,^��77�o��E_uŠ�ʨ�"	+F�yz{Rr��WJ�"��d���ut�v��	T{1�&x�����{�,1�ve�`l���yv�|(]]#��~��	�$�2�r����-7?��a1���#J�e�xGӊn�;�:]���K"]�v&^�:orOA���b��ms��P#U�Q��&�|z���+���.� ��L��o2��=���c �oZ�4Ɲ��}��ܸS 5�1	����(��}�\���^l �!�Y���X|��7\��i
�Z��)R$��O�G���"�eU���p4Ca�f2N?�<2�ͧi_�J���񉨶���Z�m߃6�A�!ǞP��vlZ7-�����Ҍ�G���@�z�3�,����(��#rp@H1���j�,p���L¾�>��6��i��.e�o�
�Ŕ��i'�u�>����@QN�s�eW(��F���G�ύ��E\��!�k�G����p��(�#p#0CI��C�Xŭ�}w8����,����>��ǠK&oS�H�iL�'�\c��wNf�H�l�J���r��D�o�\�A� �]V,�X����������9H2RR�巖#Ibn��!�#.٪�^Npeӻ/��30[�\��<Ũ��I$DH%ǭ�g�b_%[=,�'-�Y�r+T\��rЙ^�8�mp�i��3�wk��m8�DtN����¡2��*���S)d���m��d�m~�0���@��f-��򮼡2�?5��ó���C��2 o�������Z��q��*?��
�'-��$pˮK'B)YN��e���3j:��4Gs�B��}5�?��
٥�of\A�T��`�9��8E�6���_��@���Xg8v�:���}����^u����HjЌ��O��l<�]l=� D�ט�擛�Ng?�d�"�[�U�~βC���F&�g*r���Ja��VJ.x@ޝyy�td����a@ώfȻ0�J�hgc���-��.��6���i���\�X'i�I@���4%���4�vf.Y���K0���S��z�T@S�ȗ�H9`�^g���}♗�>}fX��*��(�}h,rY���s[���蘊7�������}�+3F5���1.�_�V-7�-����M�A',��ؤ���'g�_鯩Aц-��-y�q*%xQ@����X�@TGGnXMjY�0������Jzrc�U���Ɨ^�\��!^P2�KN�]L��ڸ��~�}w�s�����|F��"���ʸ/�Z@,w=?��ۣ��xՏą�Z�Z&A����Ʌ w6�d�L�@�ڑAr��\�k�����E�y�n�T�%�����Z���Y'��Q�c)^��p�s��X�_xk���;��o���dN�8�ϋ�3L^����3I�3&+��vk��'2�k��5*���~���;zO1v�r�~Y��5Qg��/�<䏍J������ϖ;���٥u\Ŝp��!dru$R�9ۡ4T��2�N�iV,-k7��ВS�~O���U����R�+�������;pV���l��Q�R0o:��>)	=��s�H�aP[&�t�������F$y���2M�5/t�zڗ�F������G����׍D�@�
����t<����^��QѤf��4�����
z]�&>�S�U
5:,TK}��� I�+�w��:%,�9�b��k3�{� g%��uX��S�c`뎵 ��@B��]��6�z�H���֑�c
R��c��zH%^��́�C4����3�%{���^,/jx�\|�-[Q��Ė=�|�SZp(g�@�#�	��R!x=8`pL]��9ew7l!q�=�$^�k ��'�L�;B��w^s	A��.��N�R��?4�I�TD��X/��MU�m1�I`|�ԷM���f_��!�xU�b����F]X�B�v&q˅m��u�g�8F�[6��g��@�����u�`�Z�;��)���X���Ȁy�NwM�Q��z��a:��qt�WPZ����9|n�(������F��i*�Y��%xn������r��ȷc��H�4h��M����GCS.8�q�q�&�9�Hh�дI�IA�:���ut�a����!��[�RքlԚ�~K�F��h��Z�T˩�5_q	�Ӱ���J�5�e���i	��n��t�g�+��y�1�N���@(������(\Q���4�4H�o�5�`�+��
?l��zB&���x�������F�/n���^e�ⵐݴ:����<l+���]�����ŋ�1��/0z
,����'��=�J�`x�r�Q�X�\�����"0�Z��[@;m�Z�C5[t��̈���\�v-���B�� ?S���8+P��}3���F���$'RS�:u1��O�Y������rc�6� :gA5�A��&�9�hQ�����9P��}Z)����)!���=kF��*���#���νD�~���MxB6A��,�����K �rr⼵	��)5�]�Xt<��IV�.@..�^�7��~z%�	��,���m�/����=*	{G�3�.dqZdK_!I���QBǩ�¢4�yG����f`ɳJ����2�ǟ)��sb �u��H��@��6�\gTݾ��σ�o�Mݓᗮ)��t�;U`�}<��I����8�S�o�"�;(9^��\��"�yY��Am1D�69��� �i#�/0��(����ʒ�Π�ɝ�[B�%���d0��{�u1����qИ-D�
�x����^wPe�g3)��Q����2��P���{��r��kHU�R�k����[*ИŢ<�n5�w��M��ے0��`Տ�����e�*�_�����&���K��vvΪ�y�����H�,�����G�����!���c�yw��KU@�_n�UoqW������i�FH�i���	�D�6V��ڽ�4��8�T<k�ls-�o�H�� 9\���w��[�t'�|��0���m/�]���y�sl��~p8�n�6�����I�B9��=�X&�^����8�q��ݞ��'h���^T]����{��LӞpo�7���A�r��&�K�����d��t8U�s��5�S���Ϻ�W�!w�Y�\g�üɊM�z6Z��[�.gSh�J<��4=nw=�փ��`e���bEJݵбJ�=�ˮ� �?�I!��������ƫ�f(�@=(���:��ql���7�L`�~�èϸiQb�M������7/�
�E� v�������ǫ6��}���>v��b����y�~R�7�.H�E%���B��S��QQ�O�87<�,��o�A��� �'a�´<Qn=gAr�y?z���{�*z�cŹ��X�pF&���(0���r����	!&KE��TDO�
ꭋ�A5�L���\��:cU2�QB?W3�`�l�XL��6��f�?1�������JfЬ1�ֵ���:)h�¢<%ks�CL�z����@�X:.���|r8ڏ�"ʜ�D~����i��v��u��L%���·�2{ë��s����4r�h�%]r��
��X�飞z7f�����7݁^$2.����Ѫ�5v]�ZB��)�:TZ��6!�*���\�Ll��$I�0¶�}�p�Ubt�p	;8��#�U���Y+��"�<x����z�^��60��������� "�8�0
U�dq�kMѫM�yE$�?W�im�F��J+u�A�$Q5�Zb��7�c�Äw�U���A��띶8�^n�����<�)�y����!�mВ�j{����q�75��"��7��g��2V	�k�ChY�4��s[s�yW��a�6 ��k����N%��[�h����Y�d!���D�hǯ�JI� ;�x��	��Jgѷ�%����f�02~d���Ѽ��i��΂�ܗZb�zLr�\x�j�iN�Ά�f�3K������9�e�vr��(��X�Nϐ�K����e�|AB�y53M��mkš�:���B��?��VQ�N�,o���>��2��џ���g�p	�8�&��w�������QSڟ����	���=�ݚ�m)r�pw��KOa���Aw>��P�F�������3 :��e���_:)���B��E4~(��uX�#�4nA���r�;7n�%�)H�̉�`����Z�S$Gp�f=:C�;�SoҠ����>�}l�)���p�us�,�9���Q _B��=>�t�F������$��>6�}����=ݹ�v���=mV=(��E&���1W���+C��XHQYx��O�	ؼxQrү��!��G{�1�	6���0d���G��V�0?a��x���cn�9+����ϭM3o�V��o�Xm���f�}�I�ַeB��L����n��h�1h|��8�R��
�~�CPFB�����*�� ����|0�r&;�*�
�������+���t,�vx��o��,Q̔��wBIA��ι=-M�����X�p���zf�+�{ǟ�	���M-X^�쓁m �k_�5-��	�3U�Y��v�bX��L�;�R��'�����\���U_$r�!V���i�g���L�)Q`Hh&���������J�Pc�N!)�H1�
�E�i�.���F��1��#�N���,J�B �f9+�r��A`�@);��9�g����֣}ZP�bMl\��Ӭ6\Z�d]1'�(4yc��6Q��!AN�G� y\�]:�53�CM((FUl��Xo�ՠ��R��tb�-=_+4SP˶�Ibw���� �V����q>�03�{?o?z�:'\tYP�锬��{c��'1�c,��8��#�I �9>[⚛ж4G��:]�Ke}����u���0x͞�~�qC��B��mn7p.1���d��0��>P�c�z��5n?�����,0<GP�~�c�u��ȄB��J��;��2�n����f._����K�0B_���..��a�;��J��j��~���V��
ύl�,�ۄA�4,���Z'x��3gs��GV���� ��j����Wj�?'2�;˰��O�2Fi���7^P���k��J�] �_��tm�4�d�5�Qsg���h�YP'a�p� ������?}�dXf��M���Y��%�1I���^�R�s�ﶨ��3��ef�軑�A�^���l<([�'�4� �P@�v��b%��ja��E����������cw̺��!I�ۂO�%N̎�M�|���%6��[m��;	�Is�R�L
���F�p��㙤�[��`�#Ɵ>)k��3qU��*������Y$��6�˿ć�jY/d�1ϙB\�f�C�F�J-�X齑m��9��?7