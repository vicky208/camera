��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:���[�Sػ͝�MW�K~.2*�����;�+�K\"��2�4�Y����xl�7���JM-Ư�@�q��>V�w+
��g�������64�'P��,�����:���B�����5�%j&Lc�:w����)�D�qR�!�	�u�A?g�m�ϭ�MA.q�TTX����%1����P�P ��S�@`!�D�-�E#/�?�Lm��:;Y��z@ƚ��L��קU���
"�!y����[�r�T]a�;fBY7�9�-ڔM�A�y�p}s�E���~��S� �OL��+ͺY!a�C��!'(o�M�W� �A��p���o��{ο��%��&�E���O�C-�.���l`��g����W�2��1��дM�V	D5g�9ʁ"8_�_�qV��Y�Ou���&�1,��Z��YU%j2�Ѥ�R���9oM�۸�Or��K�CUT(��qԌ�d��I_�+�Wx�3��]�V򥈪�S��k�5oXn�G�۩jSSy���ܱ\��c���{�$��)�R�4�6��f�V��L����QčS⶞�l����nϥ��ڃ��]ex�9�G�f�a/@�&�� ��p�Ԫu1Z�I���+�NK���o�T����d%O��I��f�w���M�4n,�m��Ey>ԙf�{6�������ՆS���<	Yxh�{c�F nZ�T��Ѡ��x����R`��^z	,=�,K`VD�-��,��=C�W:}g��:���H�ܡt*����-͟���.e$�`P�����ZZ��P��\Ȗl����pIo��پ\H���Z�B��Z��R���~�^|n%6/����ڒ8o>�ߤLT+��a�誳�����{�߱P�ڠ~�~���Af�"ckޝ���"��=�ASB���M㦬H��ï�h�Xp�;AH��͇kq��X�z}er��Ư�W%����w|a�^7�S�P#RO_{��k�I,��A�;��c^��.�a����p9�^��/L���9c�,��E2V���G{3���ۡ�r�BaP�m�q�k�[j.֗�:��cc#E�Px�a��X�Z��H�^K��+0���~i0R�j�j@�l ��Ʌ��O�׉�bE
'�D��J�����K~�_�#u}������� �l�R;vYEh��'����zQ�x�n�)!�K�g<[n��KȀ:���%�����N3����9l�7�(a�M�N8p�.�	/����f��Z`.
��>�a�/{�N��t6~ˊ��D�%�5���8v0�>���sr6�R��ˉ���Hd���R},�0[q�,.`'���2�*�l���?j�w��O���5Kg��;X�	M��am��@o��rǖ��:�a��jω>��s�!���ʼ:��ˑ�B��0-��>,�o�쿍O5�u�yO(��m>U��rӝ�X�G�m��u�����V���^urA����l/>��q��u��Z���Jg������=��e����7sn�|<�&TUI�:�������A�V��=�#y4�mcQk��l���(F%eS�ъP>�QAh@I�G�}�L��7V���,��!z0��m_AL�؈J~�ˆ�G�3�����g"�����~��U[f�%1"0�w�����@x��t������!Z��g����j��7Hk�~z�㷪ؓʄ:��T7��l�K��3�K�?�8��e����1�?w�A/���e�Y���- ���]]�n��ʐ`���0�b�;�9l�,����V9)M翆�Z}i8�>-���Q,���A���A��񓭭H�- �3��_}��M4�&U���swѸ:�� ���h�Oc��'߂S�Å��ZjvK�Իzv�8�v�\�&XJ���~ѿ�TӍ����X�=�ca�`���Tc7�%���M�U�� ��D��*EuA}Kix,m����FG"�fg��>����a��V/��p���p�!3rJ㪃����GT���g��4���l-���u)����s]5٘�k�j�
Ά������^��1�e>�EY������Q�)��*��+��!�[]�~*}1�)Rr��b�e��?IF��� f�����EP8��5=qŃ�|��Ԍ*�8h,�>�
P`�Ƅ�[��{c��Q�'�itX{��~�ɠ���x�;lb/���e�:�z#�!�`	P�����#�yw�	������MdX�ŷ�I�����DX���0�*��2���,��,!��
rЛ����e�C$��2@���8c�C�!G��>|�4����g���/��M�X�t�d�qAA�b\l��㿔�����Z�B<��d�c��1�y*L	gӿ��-�|l��4.�X[����xjES�r~��w
���6�xz�Dn��K�q�wl߳FK�ֈ��>��T��7��e�8Y,�N��?��NH i�Q�Y:>0V|0.A��2���ʃ:a��߻>�P��#�xғ���0^��[~��\�"��2���<��%�AݗI�?�}]a3�D����&�n���G���K*x@�IJ��IS��"f�03h\���=ky�nr��[�F��2n�KQZ���� ���)�y&���|�
pJ�ֺ�$�|���`n�ߦ�S��C��C�U���yߝ^!���z�i.5n��ϲ	��	���ا���+���q\��l�kb'�G�۔P=((�2Mm�:�������˺�P��X����������0��a�����0�#N�Ͷ7���o�4C��
�1"�έ�_�����	 �c����2N�v���+}�&�YB#����"��w�9jhF`�K����=���7�&���-���H�ӯ[���!�bs�&P�,�����X��Mu��I�:�gzDJ��EA��x�D�v~��u�x<Y�%G>��w��$w1�ī����'ڭ6�3Jv����yF$bJ��GNg�uB%RX��$��%
�`dĤlv%�/�Zz���M�}�4��H�Kߛ�M�AP�b���((�%���	b�?���^��T�p%�������1�x�`y��$֏�پ�utұWU�Tb/���,�/�n>E��C�C�Ji��K����֌�
J��d_hn���{ʾЍ�m�X-F�V�3��`;j�wὉ��*T[S���S��X��!fK2�������q��}\Uo�%�OV��׎�)4�A���h�,����[Y�l&�2W�G�M�H"gT"��]C��rcԹz�G�fo��6�a��X��0ߡ��Gexre!�9 2�.���l���xkq~��ډ��Xe���{[��}�B{�g���Tt`>aP>�\n�	<�`d����W៾��U��Kcˀ�x'���N�:���$��D\��WW�Y��-=����ݩ�����D��N�*�.���n�P����r"��汈� �L�#!����2܎@槆 &�� �y"��gQ��[)IF��B<�^�█r^���� kT��\�XZ��I��G j��Q�4W&����� �*'+n�ó�������)��5�y�g vP����gpN�T�#�1��������[��m�!t�E/���4BY���_Ϋ�/���t�`y�i�@�s�eƣ1�Z�Of���D���h_�6����MI��G����0�d�cFŐ��S��^g��6u�)`*����4�'���{�Zt&�?Z��s����Q����<is�̘������c�G.g	�x�='��>&D�K�ܗ&�N�#̤0�8C��~�MO�4��eFbg0��ba$P��H��M�gf��ƢO��ݰ-�+PІ�(b�p��D+61B+��!�y?������NnE�9��ԏ�� �n�m%�mfw���9O�4����b1��^�W��L�@�rmyIyjKx�Ȼ�.�d�{V�ս_�����R��)yl���D]u�,��ː�����p->X4[7=4Q�]X3�m-qt�e��F��kX
�Ֆk�>w�� ��/�=$�A������@�G_!�Џ��#`���[s@L���s(. �t���U�>���`���dQ��\�բ�·�*-5:Ɠ�Ap�\�ݳd!dC�{��� DП�Z[Z!��o�PP����/��t�`�˷��ʻ(ݎT�m0�U���Q� yd��迾�(;�C�r ��>�	�����3�_PA�Og����&�B�a`�ϡ� \8R��V�6�k�����>�ۓ��� �u�k8�jc��̂��;�^�� ����-�� 5ξdZV��:�a!�DƆ�G�k�h�ձH��f�o��k��s��w��S����9H޴��I��)1�����&7�QE𭤾]T�\�[Go�HS�A@�+X��5xMf��x��5p��p0֘�R(?�S��d�yϐ��u��e�LÎb��%���l�^36�Nq��ouF�,�~/�e��.�?�>ߢ�;����8]q�U:�U�3�4�rT�ʒI���e���#�����(?
V�L�D���iQ�w�Q��{_�k���S%�9���I��H�-���RcO>�3����'}�W���,Nn+���٧0|ZD���w=������0����G�0�!����k.���{��K�vT8�o+g\���g;G'�Pܾ#��a5͊���xh����'���e�㞻�13)+��JT%��`t
���.�g�1r����vv������Ed��H�zQח
>�����顇���?cK�Ҥ�����pˣ$i�*e��ߥ����U���3a��Į}��� ���M�z�¦�n�����~�9��*]\L; +�&�q�	��ST���b�*ի[�j=���:�)e�l�����8�8ZD���@�m�����(�	���W��Ђ%���Z��RE�T�����2m����'n`AID�.��xa'�b����:�B-���i M	K��*`��(VeP5nx!uI�T��`�w)�'��nl�.���K$z�+��O�f�� V�R����L0*�����=q�S_b�<���8�����n42/n�d��n��{�K��	mo��z.���7Y�U��@������Pռ��N�Z�w��p���lh!��z_Cb���8<B~���?j�4���U]÷�"�s�W�R��XO����!H ֻj���7��\tJ��L��5�����`�7?ʞ�?g����ab��p�w�L��l6|�鄌WKp���a�߲.�i4�H��g���R��t��BJ�ɫ�V��е�}��[~�����*�MB?e����~[ެ e���p�j�}A��:2��o��\��W�P5fA�t��Zf�:��M�C�v�q�4���}I��L�ԉ@A�Z�ɜ��3��#�Xg9�Mo��Ry�_��=
>�"�j��Zeb����=M�^��[H:m�y�����k�����c 75���Ⱥ��`@QJ:2��N�16���ϒ��� �B��浴:�*�6~��b|�[�GldV��>��Ee�'�����S���_t~@��4��,�\\�2�P�
�4��p�ߐ���T��O��x�=���&�._�F�as1D�����լ�O�R-Ա���6�Uv�]��l�#y����63
����i�Q%���?	P�1ʿs
7�SaTb�f;8Dg_w�����`o�e����Qk=�)-k����q�6a�8r"�)��0Y�V:hQki��.���h�S���u�m�ROjH�n`aַYG��Q��:���Ş(�t�N�����]�=���b����ÉTx�F6=ެ��8��+�;�PE�Ò��x�è���tv�)J�0�Ӫ�h�j��E�V�eb3U�Id�iw��g�T�DF�Q�M�E���cAd��NT;3ա�*�x&_���m��J� �y��}�x�NS
tGn>��٠�[��a�����BtA��:�����3�k��(r��e�s��^������Q]-�?�[��\z@80���m}��ep��	� m*ALL�"�y���������p�ē8Q�=����y0��op�zG�@9_�Y=�i�b�]A:��%O6��6��;;���C|���W܈ٛ�9�<�2;$7MCʛD��
�:�t�I�	��8c��q�8�b3f�� � �=�Ȝ��jp��Ìuշ��(��8i�g��Z���G�&h?��y��<���i�G>U�U�'�⬞������_��C0�0�U�F�Na�H7so�}Gu��G[�D�F�d�M އ��/����߬�]'}Qo��e�T�Sw�\/�/�p$��Y!��D�8[��i����ץ�]"�6��&�x�����H���J8V㶘�B�,�Չ�x���J�k��%m��0���	2�4���̋^ =F�|ae�P$����בt��jf�p��H�f%��w<?��4��h1����6@�$p������w�}$�FJA����.I7L���v����������G�دO��]���i�;!�臔�2�V@FI*r�͔�B�2����Bj��i�^��]I�
?�z�,b�h�[:hM�K&d��JV)Ȏ��)��F�\���B_��a��.D����3�<X��M�|�W�+�����OC���O�2n�3�}��O���[��^#pa�Ao����LzD?E�F��W�A�Ǎ֙��خ�Lv�����S�ƨ��p.4
�'5�;�X�(lj����1i9��.S������XUK'��%��?�,9u+Q5;F2sgT��<YꠊYT�����	��Y��<��⋱砀��l�<�ݧ����9��4J	�����5��J=�g�r.l�T�VIWt�Z�ea��l2@��ئ_(<��n��'�K�i=�����4Z4�&$���������ڽ�ɽ��Y�L��f���D�H�j�^���J�5b2ߡ+PΌ>A�Y'[�s�)���8w�%H/e��%�L���������@�����B=Z1�A�#e��g�셓�ӂ��i׊�+T�L�����?쥨�{��G₩*gb�}a4�f��)�I����C����$�#�ze�
�Ƽ���f:��֡��ŝ\?;|�e��=�1��~|�f�a,�)4L��LqI6�H���x.�V�|�LS�Nި2kL�ў_%њd��C�8��2��;�Rh�Rq�1�SI>�nۍB�ıލ���j;E;��EQ˗ٵ_�xQ����(��-���W��`�'.l��AG��r+�.a��L]�|���dAj?�/�~bA���*�p��&�D�v�P���q6܃@%���uW�}^���*�Pb��$�k�|LĀ/���nVL�W�jM{X���c�Z���A6���nR��D5��k��]c���YP�_s�$_��i�n�����2��J�{Mr���W=VF��`%j��me���|���vO<�.��XV�1:d��QگL݆{B��Ƀ-�>Y�XC"��?CZc��-p삃2���R�N�C���7_��c]�&���Bj��g<~���Ɋ�[�J�<1z�I�-+u�Y%�o>ة��xi����*x*7��d��BHE�M�)�o�i��XƂ��TY+�o�}*���I��������H����|.�wM��v<���q@ɏ��hf�gT�7�)��>qm�7�4/�G`�-}6��@�)��cfT!�i�o&�^@)��=���e�
~@�xpQW��+�뇘K��о8��ǹƍ~���hQ��Z�o7���Z����K�pC�N��ms��نc�υi}i�e�f�����*���5�Ѭ��+%�@��NE�Q,x�?Q<l<�B/U���a=d�Z,'|��UU�kۿ�3�E�vaw%"`��M3�}�o�+a�P%��갣,�a�2��9���&.�ex�zY�d�����:�q��ח���BEDߒzv]D�x-��t�m��o��������l�䈀�|���������vᕑy&?>�卫�~_	�K
9�$Z��������H�`p�fi��-R�Bg�<�3�*��%AL����ȑtݓK7��� �����d��;|k�s�̵7��/���t�B1{�Pyp7E�pJ�5���O���^�.��r)	������'Hl\��&�%����U��^��Z�O'l�0�N���V\;�ЬCZ�=0-�R�[4��(qx� ;�"���?!!��nu�;�ہK:������W,�Y���\�Vy����p�h����,
d�*���Q�2�I�����MO=A�b�O��m���}V�YᯫZ��z?��{��)O3;3\�!����dBYzJ'�v��\%}fȩ��E��CØȘ\�������s����ZN=���)��$j��@�,�\	�-�B�zX��������K��j۬�}g�~��
?��=υ_{�Jz�?Q�֦W�k�p�F�����g�q���`[}j�OK��c�G��^<ʳ��Qc�Ys��3u��'-um�2�����T��?���v�G�a���~��c�̢efCJ�c֝����#���J���B�X�C���8�/������IWB6�9o��=��P�nɆ(&�5�Ǳ�Ќ<+���sC�Y&3=4�)9�ĝi@��vâ�FO"r6�9+c���rO4�Ԗ&Yu۱Z�Q�hֳS�|��x)^6���!^��H����т��h+
��!�'G�^�-g��nY�Z/x��G��W��{�wK�y
�A�Q� �5�\=�K���A��% �Z��o���@E����aG-y�$Hq�X�:u���.�������@�tJ��{��!��0��A�?��\+a9@u�I� ��ķrZ��	���,Pv�b�F���~(݇���4f������sZF���3.=����<I��m�^&`�?w[9&��,eQ���#j��`ѭ_Q!�H2��(j��硍�sȖ:���#�L�(������y��C
�S,�Hy����E*1�?��:ZaG��:@�*Ƹ�ּ�?�����&Ej��G�4�a޷��[���ٍ}Fc:ZZi���_�W���4��^������a菛	���{��q�<QM|��W�60%0��/;��R�9h|Ag������ع�*�@T5��Pܢ��l��Rs[y���4�/'��h8D�A�X2Α9���u���B��׋� ��u�$��ﰩNx�������l�?��h���Oh#��
�m'����I+j{���ڀQ�e%p>+�|�#SG�Ʒ��P�=z�ytI���n�f��f��8��D�u�ؔ�7:�`�GĐ�p�W���Yj��^5�y�W}�p}S{;��=Zz�K� ���@P{O��L���H�ؾ�M��\���'b���N|Ph��:�Sp�Nil�32ſ�u����ׄ�\���-����o$��ҧI&���bx��cڟ�.7����<*�l�L�e��F4�f6�%���ׯ�6�ܵΎ �9M}���h����%�β{�����Xic�k���JD��<����
��F�� 9�f֧~���tJ��.��
3����nha���U�)!W���>j��x��^)(��FW�Bl.|~Vd�?i��,��7V}���8>u=�5-��@����/39�#�$�й%�\wT���D���=��~������2[�p��6���+���!�k}���p1? ߗ���Dd��9�ȳ-
�M�g»���=�����\M"�~UӂD�s����C�k�ہ��}A.��C�:��Uyn9�=FCY��I��fxI��4�c^+*�hl�y�#pa�}�����k��]������=���u��⳩x��VmĄ��O�s��I'h-�J�5R2�kJ���'n&�}�f��V�<�z��ӑ^T��!�|<�b�@����b�XE�ۡ���?�iRq:��ݡ���Y��S���ӫ�=D��d���n�����0Zr�	��W����0��������7	Fv�L�m�.%>ǩ�-h!|��z͗u�4��/��L�Q�<���O�P�	Ǆp�W�YX���qNf�P��� �M�#O�c&}��B���*�'��\t���-?Um�O�1$J̨L�;I�~����/ȟ��!�2,8�Ң�����pY!�Վz��Go
Ë��-V5��3,��	4����\��������W��4rB�ƅ\�����/ؒ��t�� ���e7t�?�5��tn�0�Iev����YL�o�5l1��8�	[ǌX��B{��>�ԂL�����:�l�֚��Z59��@J��PY�W��k(Q�̠'R���뒦������aQ|8G��#_jY� �ϫ��'�M�pƉ�A��EwO�L>� !QC�����=��gl��N��>g���������=ڈ(�f�z[��+H<�{!^�D������FY�z��B�7�	��p��K�	�4;��dؠO-��݁��tډ�ܒ
��P�N�n@y�A	_T�Ա�����.��&վ�:��Pᥥ#\��[1���bL���=wZ��C���^'�K���m���߾��<��	a�/A��������.4BZ2>@h'Y�nH|��T����J�����nH3˞[��P�;a�"������S�t�_�ߟr&�W��dr�#�P"�Đ�.><ɮ������&�U=�/�Ӗ�T�Օ��H=`���:쨌�*�/�-'ֱ�zƀ
W-�(�� ���h"�R:���g2!Ӝ_�l]vG�s��Z��SUM��(f��*��q��DxF��o���s9�xn�b�~�k̤�Q�6C�qsDH����Z�b(=-0�#��C9��Xm�h9Tr���9A��SR��(s�4L`Y#�K7��6�n�~���͗*4͐ �zpƤ��oM�R�0
�}9�C7��x�zg�Y��B�ni\�2�ħ*0���7g�5��l��r�+◤+/Ї.w����N"�h���|�_s���,�q����S�e.r���䖦��##����� ؜��?����+��&��>��Oag7���Ͼ�����v]t8<���<���J7|�N�w_T�Gؙ�_�dI��)�Sн����b��I�]�O��.�}R��N��׊�����3��ӧ�q�����P�Il�2Q�"Zo.5�C����JQ����?��|��"��Ri�+�2Z�-O�v��ZVNB�?�dzY���N��xd[�/!>�܊ug�0!x-
�K�O�_5s�R���J�	�}�c4<���cԎxSb:��S~�?���χ�5�ғ��3���;z�-��,�P܀��Nt��U<�vD_��[��!l�'<|�⭷����$��C�TT�ܞ�Õ�� ���-��H�E�4w]�z�E���}-@2��f�*9�'5�7)w�ơo(�~Xl�y �N��xFǘ�����I��f_�S���>�Ep��[b�2�G F�W*c2�=�tXV/�o̴;�{dTXiO�[��E�ӱx˃f+-pT��0,"/��?Y]�a�!}0�M�h~J�ь1g�G��;ca�~7$���*0d�WY��0��d��Ϝ#�k���`�3`LI8�dj8�k�[�ri��Gkp46���z���!(Ћ�����V]z��@��S��.,��$��ؠ�0��.��J�ܧ-7O�_��F��Oq�-�����?n�F�B�FH����R�т��2���F�$�	�x9���S�	uך��^�,�N��o+�U������������������"
�_�#fv�R�
�^<�G����
��b<�7�r�9�5Z_mk�+�
ts�v������M�'$���o������H��6#lG����2�
<T��ӻ��3̮�gK2�/S+[��M����X���{E���߾��׊�� �!_#��΃e\R�g�զ��u�T�0�fч�o�
���,�j ����j�|tC��+���YgZ��-�Q��Ȕt[���lܯ$��%:F�<����y	.�`E��9�U���n�?T�e[�ޙ��2%�9+E{�UT���:�D3!:�8Y��T�B���a0���@�&(rE�Sf�$����k�Y��"N0ya'�c�Q�"�^H�e�3o����3}���k%�h�[17yw��43�@CW@{�����`�dʟ��]l���
��t0+W�Ջ ��4;�į+=����e0�P��bÆ�0��`���P?3;��|�Tfj���^��c,��l2��+�/���O����h��7 �����6��s����,��W�4]�GfW���=��&ŭ�}I!���9�p�&�i��Q�m�Q��id"w��h��=��h��t��X�+��Y�S����8 �>��͖�:ܓ��t�(z�GX`#ݮ
08��v��*�j^�vq;�]����*x�cIȳ���~7�f�tD���Ps=���Fu7=y �;��w�;ę�]aN������g߶�qᗥ_���zȺ����b��һQ7��RN�SXZ���K�����~��k3���85�U��C&щ�]�W�R�pw��Y#+0�]0�+k��m�B�v��O��BY}��E"���*�q�Ǧ�	�t�A?�c���͆��(��u_�T�Hƌ�� �p-ۖ{|�ʗɅ��j'��c���6�y��g؆��ni���h8;�>��R�\���YK�R)�&69��xypB��Vun�.e�̽��;�ȁ� �Ҳö�4r�0�%�������>��[�J��RU^���5�i�U�74Ìi?��j�B�H[��� ���o	��փ�auJH!\8r�	*K����G�>Dĵb�����,�I��/�	�I�K����	��W��	�1/�&<���r k5*�R��M뗄������Xo��eƒ4-@L���6)6��ϙ�d	ፔ���G3��;�5������)H;��j�G�هׇvȳ�'&ה�W��S�˧�-<]4�z2sLD�M�	��wR��p�	B--1C	�ƨ����"�CQ��^�(c��	�(���>��Sd��f�S"�y�z�;*Q����h���Y'���W���9�b�������~�#K'Pka_�3���6'}����E��$a�u}�7�f���I�'�D��E��!
(�����������r��y�_I�e���K��<�it~���85<�@�A��cT9t.���%X>��/4X��^_��c�X�;�YJ�tN�Tz��'>�o/��w������x!ސ������΅�-�@�I�1�iz5��oh�p��I�[xݽ���D6z�<��LJ_r�^�_r�|��/Ӵ{����X�6qa	l%SҗT��z�T��O�w�OA>b�B!��V��?�������B��$A��p����w�:Я��ܓtEA�xe�~)�}�5�D嘽���,H3� ��0_j�ь6�1U�哼i�����8�E`�L/"��>	�@��ɡ/~�x��]u��H]�n��%����0�Q܆����6���~����?����)�B���P:I���ٙ(l�d�Ng����t�bƀD�
��q}D�?1�0�WȐ?E��ד��c��N���~�+�׿��k�'�1��SVJ�U�bl�������F�2�x�FQ�Hz��s�;�a�G^ȓZ��i|���p�����MR�v!�ڱ6{��W����7��f�=� �q�Cj�[���C�n'.�Ms�hX'���'�g�@#,f�J����T�OJ_�, mН�K����a<ޞ�=�k�/���}i6([E�'^r}P繤�7�z�p��Pti)gB���݂"�-�:����E��ZW	ly�ڇQwZ�D�8��YB�Y�#I�-q6����F�~���IA:�Y�(v`�{n!�=7�
Bu�A����B�v��#�֢���^G�"*6f.�/{�g���
��&y
�S;X����3)���%��c�S��\ ���4�HJ���/zz�
����J>v�>�t!��{Q�6��/Vh,�(��	Kϡ�33�ϒ�܍ڤ\q/]��m���}������j�y� Z�k���/�G-g�mw܄�AK@��-��:z�F�K��O����&sޕB5ϥ�1QEr~�FAA�f:������k�]�:sЍ�E����v0��:��n�W��~5
R�ĭ3å�� ;����PN �=K���n��lX���&�pړ����*��`Z��͋;Xm���v�/�"�JM	�H�Hy@��T�Q*�G<�@5`:k��A�q|�^/(����{�R(-��H�LY��_}��>�s��T�J& �o���7�(���utS���VQ����pg\<����#�!����rG\�̳�5_{�[T;�dI�x8
�57��y�`��-�]��o����B��:���?س��5>q0R��@����}�]m��Sٵ�F/:N��)2e�#2�Z���*x�[Ve>*���;�K]aKҠ����턙��%�鷹E��?R��dE�Z}���P
X�����=�h��
�s����x��:������g^Q)��`�+B�cJԘ]���B���	H/v�����Fl~�+Zx��+�I�|�˪@�I��>�Z��UY�\8�5�ϳ�E����`��H������K��.l�"K۽�H���k���c
�����{���C������r
l~�g�,�r<oTū�o�u��w�	 _?l�xⶺ�K	"���: G|w�ڄE��
Z����b�����]��F�`������1��6v���L?�ǈy^�k�m��Ӛ�,U`�G���F	N2O�	."��XG���h��� w'��U��~��nÝ%e�5�oL��t��T�V��B�����S��?;Λ�G�Ԝ��K�0��uRƴE�H*+W>�	n%?�D3�I��&����kh����t�7�ڐ#t��s:O���k>����e�e��)�қ�u L�ҋ7)� �S7f�[�p%��V�mR�y�U	��� l��⋇ղ�ժd*b���l�άf���mA��.L��԰��_��F~��WU9�?=�����c��<�PI�f�C�Ы�i�/ض��|����	��5�=�K=��"�����������e1}.;Rj�ƙ]�ђ ��=Е��^��*	�O����m>1����&!��J������F����"8L�\ ������W"��v6�����?c��-*SJ���>�[d@Fh��$c�U�;ĭ��(�>v��ߏ��K/�.?	�]��&��k�l���b�ԙ,p�;�����H��'X��"�?7);���t�A1L��[UкG�����̷�K=Ő�,�!� ����IB
}X��8-�g���)��Vi�����Vc��iy��VTz���tW��T�@8�H�Ѵ�(���T>c�G�K-Y�Wn��-o�m�v--U�3-W�i6��r#�i����c���<��{������AO ��꬝����#	;�_G�beG���:�P���(�\�-�� Oa�Q�Z���F��y�U�>ޙ��;1$����şC���6m���c�(��q����u�?p<����'o�)LI�Q$��a���k'M(h,��7����L�uڥ.�o�`G-�51ւ��C�ޗ���k.�b�9����Oa�ݝ�|���Y��ã����4�2�sl�K�i�)�95�/�P�BsE�ʴ5�вs���S��r$��w�`e��H��D0�n�QnW���+7t���Рt�,[h�%x�����X��i.E�v���(SF�ٜ(�������!0�C,���Q��4�-����7G�Z�#��:xl!�,�����|_1��b��55C� \��P���lqm�ԟ��R�E�5�PY&����sY�T�$On��h�z��{��r��P#�;=�t4����×�nQWR����1�0�mH����ūGs/�~-���A��A�z6*_j�D��w�>�͇�����u�!+�;Y:�䏍�=4�8G�5Lb��v�Kῂ�1S��7��SL�֥sM���NN-���|��0��l>ͼo��@�n�hxl��E���D\��UcU���k��c.�T�}����~�S]+_��=TL�8\��U�4U5�Fe�B�����<�3�%*�m�ۃHDJ�}ğ˂(1��G�P�Q��w3ՠ*���!�ّ|�i��X�d���a��95��_�tMj��)s�|�3�v�X=Z�a%���Ǫ�$xsD�E���a/"�Ż�[[mk-t�\�����G7'��N����TH��b�������Dw82�0�X,�u���H9�2�$D_�4����J;�.)���/�2�?���I*�Ɣ�^����e���E5�eJ/YR��� �R1�S�:=>l�%���EZ�wk}�"ֺ V9W�X�+	b��K,]�.�������,�nx�K�h	-�+唲��-�l[�:����7j~p��v�	�:�T!��I<�in,"�B�$C��9��afsL�L���6�����ey�]\�4��J[OD��1n�?4۷�K�eո=33��Ψ�(���p�H)�z��Y����x�F��kf��I���{1D�Fj�4�[�P\6�b뒴b~W�^9�Y�ݦ���B�J�0����3��U�|q�n���䒶�\X2�ר��3<j��B���M�\�:���D�y��	�~[\)��[����7�N_�#fjw�y�:�u�x����
@j}W��԰���=�8Fo1����2s_!��\+lX���ş(�[�lb1�)dA^8�f��:#�v�np��KUA�>u��o�[.&'z��٘`2{��U�M|�ط�?�������,�]�V�2�,l;�M��-���lF����x��!�1���f4� �Բ�L.N!i���Ԙ���[���f9�z<r�u�B�䁪�,��G��A����r�%NȯUٮ5jz�欄+�x�D��n7�_g�Jȃ�E!��s�d'���0fK�����^�u$bܜ�0�P����Q�����C ��D��L.J���O��5~M�%6)@������x4�F��ޓko���0�A�#Xef�a�92�J*
�Be�Y9ѓ��H/�l���R�>��F�5�
��<���ja��e���]��������7�$c�Ϫ-�_n��X��  ~m4o�P?�`��(�Ӗf"�ʈ~Õ�i��%ӛl���\��Ҹ/��g{�6��o���2�)#� 3LPc_�7���$+co��JlbA����fM$�	::g$l��U��2�H;����bh���%P�C0� � %*�J�J܆�~셭{���M����!?��j!v����N��K����~��*��Q�pN�Nur�℉�ބjҍd���{�&`�Z�e<����]a>�3��J�?%f'�ƷJ7�r�ײ��t��@*ES+!+H�2��x�K���t-I	s��q�
��W!E�����G+G�����u��y�
�%��	�d��$|Tm��j�n���H��Hջ�55jW_^�_�o�������N���ؼ�����7C�ؘP���?�d0���kK�8�k�}���굑��e������ ��t1�'7+�����Z���xi�q��f6�Z%$I�/�����v
�Sֵ%���bj��6� �m�Z��Y1������o�u��I������;���-&�)��د"�`��ZY^i���5ːీ&���K���k�r���@8`�H)�7nM#�B�H�b���g����I��RTL��8=�Շ�'�&[����3���>�%vx"\�t��a`�b;�Sp�����-3�~�$,!܉�
������z이�,��.Ǘx�K~�<� �ljLI�"�hcN�S�O�s���'d6k�Iw<���[�M����
h�Rn�n	9 G�\�nCy��*A���>�<0 �w�F�;���|h��w�6Ku|�Q�\�[���Z� 3pz�`M1�.T�yR�V:�τ���-�v$��L�ܧKbd���Q��2���g���o�8� ���k��������I-�9'9H��È�W� ������#?�Ej��T�u�8�'�	r���H��֔�5v՟r�	9�*h6l� k�R��a���V~w`�����x+6'������ \1�M�H�,���e&]Fњ�'=�T��$�rF�BT���#�3hīa24��� >���i���=�^$�	�b���&�t^9t�cx���zh�~_�p�d���y"cW�ƭ�:��~ښwG���Q.�o,��z*?n��r�DsD-G77|~���!�s���98�9�llÈG�{gy�7C�|�mϊh�P���ڭ������b
��ߑN��*Ԓ<��ڥf��3g�̛��-��3����gE͒�xgN��k�PH�F�?'�
-kෳ��&�5ā��7�*�%��Yl+�Ҏ��R6�J���?Ƃ�������lⓩ�_xR�߽1�>�x���p۝�.p�'э *,��H(p(
�P���K3���r�\���l�w%K�̺ʯ6m�
���j�?kx>X9ڗ`��u�o^ͫ|���B�{�`��ǲ}ԛ��2m�Ģ�&+n�~�驍�����g��\a�Q(5hd>y0��B���E�������؅��)��J[n!y#��(�^�tb�����Y�/(��Ƨ;�:F�D%y��kaد�G.׫WNRﴤ
��_��4�Ͳ�4��?8�"3��v]� 0>���-������.�Yþ�M��,r�Ͱ�2��l��^h{�.񺟁���������4�ӆ�/{p�S��!x6��/#f
[
	���^�˲���
���<JF��b�bl�y������2�ϟ��jФ��;���o���e*HE��n޸�v�	x����s�"�#м�螓�����vcx
L�Yι�����(#���4M����M=̡���$A�u)�ky$rE���\��&���2wR$(pIp��*�K�����l��������~7��o�W� �̼A3=��6�raKX�O�Vn`0�zU;.v��43G�J�u�]?p֐@�9
��[�oNn��c�F����������d=r.� hϗ�ò�8������m$��7�W)�*�����u��F������l�T�n��⿤�Pur����W�W��Smu[���:��L�MH���w<�<AP6@Y�O�Ͳ�k_�~ZȎD��q=�)a���u5�z�����ev�bM,d:��l)�#ߗ��m�Ι�lD{i9��?p�^��X���J�nߝѮ���e�_̚R[:�0�0�s ��}0hKi�u&0�&�"r��v��������� �o�D�t�6��]��Q�~�������erC[��C��%�]YӾ��8$��1��K�)�%I�-gYS��i�0}��-v�c��U�YJ^U�E�!���/� ����B"BDSd�+�@���{��i��ma�VŇ�*	��)�Εm�O���.U�b�[A�Ԃ�3	�>��!�o��&}�Y9��I�<�4����nQ�6*!7:X���{�f���.�,��I>(ȮH��J_l.r��]��\��e����d� �B�xd�s����8/8�M�$�ы�h��@9�d��qp_�\,�!9�9����L�]S�f�j�!>�Lf[!M���U�kf ��3߉�sq����䤰=��Ֆ5Q3g�Zu���Q-����Z�O>DFl�]�W�K2��������0>9�r�$6��i����ͮ����1���*Ӊ7?���՝��{��M{�g6��H���5���d6�!<��Arr��Be�eQ1yd��AJ#-C<���@&]o^ވ�2Ӆax��l��O��%�UX��YK}���unJ�R�(��oX'lDz�K�<-˱��f�Z��k�#�׊�T*���mf�뜸����ٿɽ��_Kl\�W*|�Z��(�I[R��a7,t�^���ʪ��_o�8��"�(��|�h&�g�#�P'��.���C�pE�2�+N�%���A��u&��苂<��<ׂ������N�PA��D��%p�	��A�O:*1�E��$D���,.-��J��G�Uw}�
	�Up<�y��� �X�hN7qo����2ijk#�`�p��Yi�������P�$�C�h�"=_bW;����$�ˁ+������9�1���PdC�:���3r��Q
*�lg@�]�����$�4������n~���64��^���/~��TE�N�u�&<��Շ�{�AYe2����A*&��L@� @#ť=Wr��9�%<?�W��E�>�_�n{���~��Ɩl�:g��c�6u��Ֆ�j�zj���H}�W��N�c�k�0��v�|k���L� �����S4������jt��a/h~��0����m��2WNUZOJG%5���콡Ȝ ��$#!`M���:���ʶ�(�w��p� �vS!�T���qW���4X7��č�.��bb��d!6��PDέ����=h��5U;�#��p�poi����`�^g8�v�M����n�C���D�0s�U��%�h�gN3��U�c��@�3;�FN[a��҇��j����O$���5��%�/�����c��?���\�r����$'r{�_�CG�)䎤��p�u��k��/9�d�@1KN�����⢊e2��{�q��^��#N�i��#�u�0�*��̰Q����_ C�lq��tv���ץ���:ǃ���G�UT��}�����Yk�ZQ�$�����2�A7�Zt�Sx1~�O��A�c���W�����G0�4Y73���T"�+z�`ۤ�aDe֊5�i�A�5�ň=x�F�3���� �Jx�%�z\y������a=�4���c��%�zeuo^X¼QȜS�,P�۸�B���Bb�x����
JC�ӸnϬ�4�ɵ�*^���zR�,.�[�o�h~��ݡѬv4d��]+�*�H��4�`D��Y����p��[����@�����7N+�5P��y�ny-xi�� �+�-�ns!��Wp�S
���I�q��H���L�|�1�|yy��9����be*�I��4��it�6��Y)�ИR��p=�{]vE~�.��ZDA�{�����{&�J�^�8AY�z}`��
���S;�iT�4!.T�D�6��\����Fї_.ۏ��]�#TEQG$x[�e�C���v��-��v�駃�;A�~m���1ס4XȪ9n���ڝ�8��S�f|~�N���"3ؼ�1���2�y�'j�鴬��_ [
	qk09D�%N�A/N�H�Mm᠑^���"���Cc%@^��T�թ�5������ןo��֬s�Px��hB�s����cTE�yg?��?�m�j�`/�Ay��;OaN��˺�f�t[0j:�R�0~�F{��_�L���_����Uv� �r�R���dG(
Ew���|��� 6���/����q�`:Q�eTP�g��)�x��z��N����2=A��/
��:
�%�ݶp��.˨��]�7[�h+@��OA��n���SN�{�^�K���Z����@��.����k�*��ԍ?F���Lc ���Y
�y�����%�g��a_��%Zǐ�#OB&Еx^�)�o�X�&�����9<�D�R(��ŵ�^y��)���G�����'���Xwa('S*�Y�֎}OX!��x%���nș_���C/�F�~����%uoeը'yd~����ep0�\�h�:�{��Yt�K�bB�*.�T@��H���R/Y�me:�m�%-��c����QF�0:f��7���v�������D��[�ک�'��b��q$�^\bb�zD}�/�Iwa����r��#]hHw���X�şE��5s�h4�,�>�]�_�
PU��p��Z,a`mщ��.�����u��́�]�#HV�ۿ_>��Y��� �mӫ5�3�ib��H�,9�3b��h��ے%R�_��K��U'�5ŷ	ߔg�kJ��uV����VJ���G��~��?f*{�N"��$)�,�j~>�~=����XQ�J�ek�p1�$��Yt��{IJ�OS��f���񭣅�61�F���}i��L��9��Ц,�W�C%p)��z��c�g�k��*PF$��,*�����X�rnxU�"$�ʰg7� }yc�C
��^���F�:sBH?[ڏc�2�?�qS{��%�T��63�+��8C�h�q��eǛB S�0�{�.v{�4� d��6m]� ���C�*��4� Fx�����7�t̍
�?���:k����`D��k;�6~h�)�a�_/�$~|߿�	'����v�RëP���i�Q��қayY�dV!4r!���:�G.,C�����n�lUp$��������qH7�K�%ls�X#�����e�(���9�κ�����0��>A�L��xP����W�(w�C�Q��.fG�xK�]�Ս+��$���4rv�h���%���	��]阑�j���,�L/�&:�}��K�a�td$=_��Mx� �	�ik##�*��NB�Y���n�t�P��2�F�iY������;Ò�:}�W�4�s-���"�ׯ����>��%^�ڦ.N�W\R��v
�|��Ec�B�:��Tg��sYT~2:ђ\P�|��jJ�B����X�bo4~9y}.��X*QM�)K��>����H"��'` Ӑ��q�h*4T�E�W@���︐O�\F���c�Vm�z��b��U�R7d��E*}��y�C��� �ז������*5�M�ދ�u6�E�Zw��Z��-��u���"��wa�`���Y�q���BΟ7��U�,Tģ����JANXuQ-��Dh}�'��>#?��y�<��]KT9 �LUJ$	��OU\�s䭢Yg�R/z3.���vo�iD�'CI�`����.�*�1�%�7�$������]`�4��/U�Lq_�.�מ�U��q~zP�܋ns�x `���ɶ[N-��J�*����Wc}?��ps>�F����������ɑy\o��.W��HI��c �H@U	�������s�5P���Y]�����X��T~gf3H5RX��O��|�J�Xs?�
���)e�a	��g�R���5"�4"�3��:�����ʺn�u�_;�p��쪭��к&c����Y��
O���pD�s�b�Ph3���hwȧZ��6�YТm��w���à"�	����Y:FTw���=|�c�O�uO@����RK2a�����w�;s��f/�Y�Isʠ��� A���u�����^@�cs9��y/�\�<���Է��P4}����?�1��'����|�v���KFjk
�b��M �s������8׏�s���qpmM���&nH3���>��&y�}�G�XS��7��X�om�$�i���X������D����;��K�ey�c%6+�;%F�����>��㼇�H�P�.wAE��MP\ ���=�y�<�JO�U�sp5'����q$�;٦���b���]}�^%��t^�a׆4P�:ݖ���	�G�-Ė��N�czDy��'Fg�oͰ�m%�q�$���ؓ:��9�VÇz4��O��_�R��C�RhEX�M$�
ټ7X�,#a�_�i_��.���4.�8����p�ƍ�69�d1����h���u�FCq�{ې�����,w?����V���#[�u'Һ�C�.�a%<�hb &p����m��šnr�K5�M����ӷR��ΨR蜲�Ō�h{,$����������V��qso�O������M�D��X��]�d�
W��uς-p����J��	�+��fE��Ut=6./3��ѵsNL�� Դ	�P��?���GC�F��K���H����+a�QY�@VA��"������Ka�������ک Q"�J�a�8a -AJ<���d9�`�x�b�!�V���ק�n���%��a�o=W⟌O�#�8�qF�|���x�~��+4�e�.��wӾ�ޔ6��ji���87ڳ��P��J�*P�o������C���*'yY�<���gG�ƯS$�����^�v��	v������-�5���Uӛ��g�ri�M�r������,	�h�;�J�${ �`x-��"��΢Т�VQn�Y��WAn�D�{�(3ޒ��k�ZKK�M��ȩ\G�x��� ��)y�Nh2�W��yZ�����Ձco�QN�Y�i�aWE�ܭ
 G�h}ѳk��]XQ��`�9CJ��K��7)��ֶ5W�)��W�^���������$h���$*�Q2�����}tr�u�Ш�qR� �\���8Ѥ�+7U�k�n�8QR�o����ي���	�b�w/H�W�\U�8֖�����W2�#n��k�,>�j�V�?Fa�"�����Cd��	����3w<s�3�3�_1Tܩ�B��T
�jf=�i�������L֙V��OIin� x���I�Y5o� �~��Z�ċ������ΎC�w��M4��r��y�2Mh��8S�3���Z��'o��>{�A|? w��\���k<J���Hvq ����E��h}2��N�H0Q�I�-��pƈ�^vB�X�}ws�;8�v:,��9�{s��������Ҥ_¼?P�/����Z�!mhy�Z��f�|q����p�c�_j9�ҙ�b->��p�=��u,�n�TL�;�Kl1a��D0��%w��Fpw��Ƿ?� �r��c����&w��cj���.sR�<*�� n~q�\��Hy�b�amp���T�fw�f�9,ԝ��?��|?r �A�;CC;�׳���zh���Xbٳ,�}/;��#:�u<��-���7.<�"zk�P�v��k���Rz81w6C�a�j��,9j�z��Uo�kwW�nh���E���8X毘�!�1��zl��S@G�U��
�A>Ck�|�9�g�W���y�h���A�I+Mx�9p�
nV��
0����<�_vo�� ��z�M�jl�S�o�,��ˋ�r ��߅c8C;��s0<���H["J2{]0,ț =��	�Ha�XY�6��H��Y��Q��CZ��J��ƺ��[w�9�I���V���K U��_J���x��x����vl��_S�ӎc�W)�c�{�r���v�i
V���^���3k�n0�~�ly��$�^����T�8�HAy���qy۔�6�'g� ��]�����0�#%͇B'̛����6�$�ڼ������)W#�����gٝ2�'�11����˵4�=��w(��{��X��8a}�,6�Yj!�bF�v2������M�]�x����AEi�'�?Pb��I{"ou��~�SW�Ul��˪U�����w1&-���cBE������X5��j��#ŒB�����z����륞x��,y���3�Q��	k�f��A�%��Wv��m�r���Q��#X����2�������+R�.h���Stҭ���v�óf�R8�PUr,�܂�j��'"�.��w
�)���f�;�ϑ�n��y��um���.�HZ�yE�����FC��׽C��L��ޕ�f�t2~�x��;�Z$rP���#�$�g�������Ճ�J���e�/ç��L̀��$PBƷ��l��͏��df���!�yP�'͟ǂB�*'?\N�Q:\V�÷M�pW%ƌ�����H`s�Z�4P����d2nEw�+����!{ &@�5�S����>�;�UAL�J��� �H��	�|Q�'�$_��a�Jp�A��T���QWm���%�k.��M�i��̱ɖ#�!�z�F��^�J�itC��?�4n�y���7�
f�/	ˡ����քjĶm���3zjhݰOP��e|H4�����������-�(+�ÀP�cY,��r]4Ǜ��sZ&�����sΣ&���<��n�̉��vSD�?c+��\�����5�I3�c�m�$pTk��؀x* �$��-��*���舚�"�q�55]O���'����
�Ԝ�3���I�@����O���&���ݖ9��K��Xu_2�m1M��5;f�'G�3(v_��^�k��S�(/��pQ�[o3�-F��z���躔��/��a6��j�����\��A�M� �U�y�0=��s6��U����#&��RD�L�Ե|7}��0��[��D�����
u�R ��'7_o���M�9U�k /�)����lV�@
en'zF�e�nT���A�뾭��x���.��	+A�'H��'�_�����}G�:pݝȟ0��� 9�{3'����J��$�9���DC��P�\V�D��Q�{c�ٷ��R#��C�/�ؗGMai��Sr����a�ݶ��{��x���&���+;�K�f/�Y.�?>�����0IS����TN� ����QT���Ql���G��� ����*����xzA2~ȺX;/2T뭏i�N�L3m߭7u��j�Ⱥ*�����h��n%�H=to��#M�N���I^赆�@R&�]��ĮVP]m+�!��߿��;�+J��]���W�cr���P��-N�MlF��XG3�[�$��[c�m�t�.�5^�#�ӕy~�On����"��G����"�󜀔��̴0�>�FTE⣃�_��g��D��ac ���`NxEy!Ce��T���9��1�j�,����P�R�����g�DI*Z�9K��y9�J�ъ�;rt����<�wg�|/k�#�7�r5��S�J�F�_�]4߆���Yh�V��':���;%��e��F��X:Mbr�����\�9�����=���:{���G���Wf��l%�0�it������5̫QQ'����(wfA�C8��
Q��4HQ���x��GO-�
�]����֣±�T;I�/�<k�"��oC�_y�.u�ۋو>(���g4��%u� �R׀:m��P�FL��'��4#3!����
h�O��Bc��:���d-�<�����S�����QB﷎!�������v��(��?�!l��@���J�z�0�,g0��D�4�˨�ZB���<����-��p�W���/&-k�r�哈�'wrJyϹ��2�b�F����m��H�c��:�*ã��������E�#;Q�K��l���Ђ�[���y����R��ho8�M���	yƭG�=�9���[Y7&"�2x(Z���W���K#��?E�+�;������'�5�����B��cl��e:j~{`s��1?���׳�N2��l{R`a��[������'�L�![n@b4�o�O=�_���6��[���
�e|�>(�4ܯ6�y����B���BM�gX���5��V�-��Cv���v�&�������ɡ8p�N�M`w��"]�w��ߎC��0n�^�4��0�����/�J�EjZ3�'�5gA��ք!LB�K� �F z9��a���N���s3(�u��j�N��<�?X=3h^������Z���!_XY3I��X��`A��E�Q i>�Өb}�ip_���w�sc��{H(yL�|Oz�g<����W�J��\_��Z����/��@��R��d���2{���큪׈qs<�+�c �e��s��7_y����I�=��f(o�w��5�V!��j���5�P�T��p�+~��k�7c���M��5p�Fj�8���C�d���Z*�(o�d=n���3�(h�K_d��:���>���rQ�eC]dP|g<@���"���5����]�a��7,N���5"�f��0j2.�Md&SQ��T�9Hx��{GGy���J�3�?���-�y��Af�{��:�E�F���{����1��sS��6zOQرO���4[��a���`Y&q�f�֠�~sg+'EN��-�m|:H����!�jd7+On�4�3��Χ�ʴ����nIw�[�Yƃ_�_��&{'�	Зӯϙ�#V7����U�T��%>�S$��,S�,�H/f�;\� ��
�X��ވ{�ײpǮ �/#|��"��
�S��(
�s���ʟp�O��7�@��} ��������`[٘J�A_��9�k��N��y"'�S�H�#�+������U�5���s��8T��&��������g�������;s}q;9�k�Ӆ����*�:V��F�Σ������6�u��e��;h�>Ho2b�i������>��q�J�	K0�w�G.2����Q�A�*�����ud@��&8�N�8����$��)v
����OqAn�Amcg��9��j�Ɂ�V�`|wf����@A4�ջk��l�)�ᇩ�=L���2$��c(��t�p-���ap��tϑH�0grw���ݯK�p{U�?~?[�v�o6�h�IxN�
��Kl���>������mf���S�B�E���6�K��pk��0�����������諍��
�e��(����HR4�����rV]G3�K�[��N�Ba&:���&p�V3���q�E�����8�˒�Y�1�����}!�"W��޶`�S+��`�i�
�b�C��h��)��K����k�4�FuЙ
r�&����9��T���!��BB�4ƿ� �I3CƋu�<�QՃ���{�ܲ������s٠����N�2�=��(���8�w�^Pw�./��E��2�B-*��"G&����O����B��I�(�� G@��]�q��ʪ剌X����ٲ�ئ�5��퓄=�)���æi���j�#/@�mIŅ�z���i�-j��X�n��	��{W�6s��O0�}Dqƚ�m@�0mWw}OS��Q9SH�L�W�ikf�/�⌹�t�8�=�@�H���6� �Sx 
�*6�}��%��n4t�c_�%k	
&��I��3H����K�3e��-���t��ݸ�"���8�A?~19�gk4��LV�l���{��Օ�"�uuPlԲ��n]S0Yvj���+)�\�Q2��z���4op}����˰��QReT���R�å�U�s~�ϛ%$��aS������ʯN���&]��BZ�|R�fɄ�*wO"�x�E3AI�&Lt��=�z��z�F:��C\�Q��Ҷ�5Xϥ��j�2?<���I��sW�*���;?%����-�+v�p�ɐ�	��>w�t%�X_��{0vC>��FmԨ/�m���d^�8��:�u}f0���O��i��c�Ɋ;u����͗�lW��(�&פؤ{���q"$����@�z��j\��xZ��P�qcW!���ǋ��UV��^),��D�"�{�����֏��+l�"JP���_OJ�5�Y6�Y���\ �x�zI1~��R\C&�2�o�%�|,ֶʽ���n����?K�(r�d;h>�Ȁ<��&|߄�KcRB��F��J���ay��?33�#�W�j���Fpz��0��;qhe_N��;�m����[�#�4�f��
�]��fgAȲ_�},�\���A7�~z��;qi���#�4 �;/4���+�P���9�FEdC�bFE`x��Hy��Ȓ'��ǖJcI&���v���f}�if�^���ߖ��p�Q�o��,�]Ӧ]�ޢ]�~G�7�B�U��b�ᅀ�ʙ�|Yq�˄�a��a�|[Z~b��b6o�a�.�~g��� ƀ�ӞWuEb���^\}Zh{�	��g��W[�j����>Op���~=�җL~ȼ�@� �	5>���g3��ϓ	�^���O�9����������O��R�Z�����8�l;l,�Bj���Կ!9 �S!q�O��ɡ�{��_���@׾�a^�X� ���%�'DOe!��*��ü��/~Q�TY����R"U/I�y�a�D�y�\�/�'�!'�jBA�f�v^e���#�
ý��^p�l��7M^����v.ʠ`�S�ñrQ~�A��T�H�J!��<�5�=:R�Y��,�Pf;�0�����=0�7�X���%�mɻ9�y��%�Q�ˣ��.�,Ǖ�+��ӱ��4e��E��$����!T#QU�S1��{d-�d�Y�ŏH!x]U�;��&�V��'<���/DmdN���_
��E;}n����3�����_CkN*��,7���A4a9�:�C��}%�=��k��+���w�'ϯDA�a��?����#�0�#`�K�����#8N�薛0p|j�LX*[��n-������D��5��	?����M<���>+�`�?r���3���"Tp ��$!3*e'���j����/����%b�����B킒�}�r�̒�Չ�h[4}��U�vJ'4�߷%�t[k_x:��r8��Jj x<G��b�x1�t�\�{�|F(��x���觜����> O*��3���]�E吪����M!jw��)��X+���o���₎�o5?D�?�-R	��\��ģ(vo#��g�����'�0h��N�)�_�5���ƈ7k4��!�8cr��u=gq[u��{D��%��A�X���^��=5}>v]���7��I��>��7�X��1S>�Z-��쌵ӻ3I��ܘ��4�,\��[��������^)�S�|�ν���'#.V푿����X�� ��p��`�$�ݥ��xKi�,��h�k�'������@TvX	�g�3��k�H;��}L�	�Ut_g9g6�U6Bj=�:���է�w�[Y�x���m������f�t�}��ժ3�av��ȫ�h�^js�E �����G0������`��v���Qm�{J9�`�pR�#5{(���0����c6;s)e>�x�Kc2
�f�l�+�7���'��ry��dd�w���A���xk�L���XC�͡%��^���D���E�E��RGVT'RT5�ә'>���:d~P׭ud�#JZ�Lƃ��z,�� r�*;�S���g�rx�?�P��g�	�7��ۭ1w��I� �n���_)ۑ���@��Q4)�:�M��9v]Z���C��CV'#�ej� �SF7����fـ�nR�ɖ�����P����K��L���� �����ވ�l��9����4�'�e1���_�y��H�o
w^������f:e���`�:E��q��Z6(e� �\�z�[eVh6��#q�V��[��so>���9Ծ����MG��/���R�����ai�4Gt%�);=Ύ��_��۹�v�Y�� ��.�&���h�eGM�^SD����+�Y�K�(4����?ʫHfk8�13E*݋��f�b� �c*D@��D���D��_�T�����w�SJC��YI'�m+�Z*�]&[&��MnF�*��p��k�·����"�:2�@s��.��r+��},W�t Y��8�P��(O-���C�U'�8x�m���nIڇj�����J=���2�>6�!Z:$���N�N:�+�hD�f|r>��L�lf��*i���AvI���ɷ�0����]���x�;�ctd�L��Q��K������,�a���v���J���N���H���V�h ��Ti8,������?�,�ۣ��*��6$�f`\�E�%�U%)뛽 ���.�L�Z!]��������?9Sf�=)FOGO~U�3|쁕��׾_pe
�:��t��mY�F�%h#���$���摬��Sq��D�#�B�A��Ʒ߷7�Y�TO���\��~�d�0v{m���.pNo�/�&լ��k�b�Zj�ަ��8�n$?4(Iў��og�'��wR���$'�g�x�CD(Ce�Z��~c��������q́S.=���x��� o�Y�]��ը��\��m