��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V�e�4�T�}`Ñ��P�F��`��^̡Zue �}���k�@��Ȩ��aF{��-&+$���������a+���J@�f� Z\C��>e]�ɉIr��=��]�{n�n�"1����:�ˠ��|�Go0e��/ٶw5=�25�V7g��LF*�>�S��! �y���<����0�K�X�� 4��|2�w� "Cɴ��ȗ}s�gUx�U^��xW��[�^��m�uh����I�kεgQK"��@�{����HT��-�8i����G�ZX'jږ��7F]/��tNP[�*������&��
*�:֌�O��1eǚ(�.��f�n���9u(���z��rFI Q{:����������
�֧�p�f-���������g��]����y��}����H��{K����/j��H����r�l�z2P�</Y��-�e�*����GL�Z���RS|{Zf�:3��{*NΈ��5v�c��}�w���[�qV�|P��0�Vu����.3���Y�'I��/��_����Y�T�4��[Q9�T�_F[�J�59��Y�1Gu@�sC�ra�}����d��
5rl�-D\��yzS�7D�vL�E����9��|©آ��� �	�{V�H-�H��ݻ�M뀽����X/j
FFl(����A�א�$��i�a�oE����%ɯK��B���T��@G|VK'�t�U�I��o����f#�񰢮r�� f��}�hL"�+���֭��o��x��:�W�� ��6y5��A��GTT�_�P��
 �߲\�����g���x+�L�|�+-y�CV�΋�(9�=.��]�#�Y$��m�D|�p���ݵD���qa�\���Nl��^�~��*%�n�c$��5��\}��d��]��:�t��	�%��F��B����w�EE���s�-j��e�	ƒ�l�<*�W�MFK�-�;�nym#-!96d��%NDb��cB��Т����I舾��u����g:��2s�C.ۓ�k���@�X��������*�����r������p
�z��X1{�~[<��V���E�����ԥn\Кa�`���]�0��[+�G�F�h��sV��!H�$��f���nbQ��Է3�[%���1��[^�W\BM�O�A9��C����o��_ ��M%�glЫ
�O/;lrģ~��5���&`W6�WBx�?��l?��!=KtE>�u�8ݬ���P9�1x���p$i�78( ����qO�,W"+u�K8�+3�g?G!x}� .�&��{Z�2E1U�_��1E������AF��>x������B�E�B��zm
�s�U���Z ����mD2h�N��0M�]F����ż®'y�W@"����=���j\��yk���+\Xx"�]#��L��q�F���b��;�b{�t�x*�MK���q�4�;�u&m�9��İ����\_��-�l>�)f�T�/�+I�2�4�+�nM�XS ��ӭ�6=�K5�97��n��5���2��_O��B5��Ʊ�|+��Z�\j4է,�"�`C�\��Tb=�>!<��Z�"-39��� �h9!O��5�ݸ�H��06v�[�ݡ��a]-��,��rME;���<ɪ[�vt 
��t|���F����2)*j��7BN����^�]qo�j,M�C�l��9�N��yMǾ21�(���$���R�1��������7�>�[֏�z33�bI�R��� 6)��L��@7
h�:%?w4<N.g^��7&û��fZ����D�NeI�@V	��T/aWmQ4\���l ]��0#�3�-�~6)��y{G�����˵*pգs���q�\?,�KX�D�
@�
(�]+�	|UK����2�W/U����W��?�
f6'^�:gk�5�Ft�a�q�Y!\8X�>`��OG��y���b�gg#o(�ҙ p|+Up(��N��>>�
	5�+謮 ��-���^d5��_�2jy�a�!���Ȑ��'�x��E3��/�O�Pp>9��i/̙#��"�U��sm���8B���=޽S$��8 ���zp�Sg��Ч�c\3W�ȱ�����k`�F���;C��ѻ*��u{ʇ_���3vZc�(Sjy,nV�#�T���؞��h4~*/C ��9�L�'��LT9��6{S��"���4�%ϊ�*��G��&��Qm8^:�=�����