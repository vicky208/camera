��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�U�v"�5���rLRU����{���8,�g�1*��)�����Vh�4���[*$�v��_Hn7��,=��R3O9��#��2@v��H�(Q����nQN�%�B�G����	.X�R��U8���@�m5��L%C���X@������l^$G��%_}1��n���qH~d1��Ȓ9�y1�J�U-���t�A��>5���_Y�+-&'�cUn�j�IO|���	@�+S��l[��L@O�I~;˄ɢ�5��q�6K�n���+����w^��`	�bs�"U<��6�����X�2�}b;gڸ���blW�~�;�t�+�'�	�z��=��31�}^M�4�)�}Q�� �� |Z�7�:1�nq�C�x�� y�=�����`��}���X�U��3K�@'�(��� 3&Z�m�/�l�h�Cm>C)�|]�Q\���h�λ�՘vbh�X[.�l~"b����d���˥馭���M)|�M�6��]�Ҁ/���Grd���m/JKt��bd��)k����(o^�Yk�22p>��v(��QB0]C�b��8_�<v�-�j?������[���G��M�����_}�~H�MY3p>t��D�M��;���VQ�	v��N�$>d� w#�|�v����v�UC/��EZ�]/�V,)捦�>X�hk����j���6��D��1�,�=7A�Maf�~�m�Ű9��8-tz�&��u��6����C�L�]�����.�U�=f� v�8�5�!�&��E�E�89Qd30�2�#]9����l��3~�9���nky�<�sXݙz���Z�L��M�`�nBWC��NI)���_m����E�0ZK̖q���RM^��%M҇"�&pf��ew@y�eaR`V$ �qz�8j��0��(QZ�D5f��<�����¯ǪPF����|����o��A��jsJ�)C�W��0�� ���:��_&� v�A�̙���L���u��G�MF������r�����8��R 
�G[�N�]�VKc��{��IO���>�C�f3?:�c�e�eR���+9�2}| B�m���Vsy�I*��F79���c��N�ߦ"�x��.ը��T�@��NQ���',�r��K��ln|��z?�"�q��$ĭ�� J�S�]��AW/h��e�I��&��"��<���ڂ��h/�2�<T��gEZ��!��
�O�$�9��d_��|�>8���#�R����3��\��{G��a K)U�����DA�J�2N�K�h#Io�"\�M�ȋ��5єS;�g�[���/�>[�W"�D�zI�.��������xs���U^�f�m�b䜨��ۓ�wh	��7
���	�z${.������5̑Vm���;��^zz����6��ؑ��V�7WF��Z�=	�����Uրr�"�5*�<�Io�:0wqń�ŋ<���]X/�\n`p�7DP��TM�=?٠׍�?�0���h9�ў��5{�6@F���.�`���XD5���c�p�ϴ\����|�L�/��<;�-i~K�"S)��L�7�c��eU��,;M�.D�!1r�<?���I�Z�jY ��GX4�xpޝД�D �P���QI�Ѝ�+�E��է�s_�2��y�2�H�+
߾�w�
8�~����=l^��i����·�����LZ�C�yVP�����w��;��gE��:�`�Ȱw@&���w��1�R7%���ll�������,�_% ]���0�]�l�,4�|�2�� �C��K)��ۙ$w�F���S�7�{��d¹�b����� Z�J��i�_Sp4�E�W�QB�J��s��7F��	&�W*$���~g�N����}l�
	xk:� ��I�gV�4�9NF�d>��+X��g�}s�+�o�u���kJ
5k�D��;83�rX���^ܬ���%e�{��s�YM?k	�X�"�)v��{J��*�#��}���� �R?�A���4s6�� �����]�v����v��\LT�w�!���tH"�s��%ZG�ȓ�d�Y�u�p�.ZǊ���(�dXDmJ�/�>�
���cM	�9�I/@����\Μ^�]�"�硴�3z��zQhVo:��ʜw��̠�9�����:���tƯ�oĀ���R�r�E�G+�Cd���y��� �;{:����ʨ�_b{o����b7�-yT����߿e攌娓I����(��2A�H������u/�nv�
��)�Qt�/�������=�*=�vF~@���P��J�["w��iэ���a�Ub�y��'�HZ��@�����/o�'���+��+K�/��� �S@gv!J�ji�lj���d��K�B��*�!��a�]���i��~-������9ܒz�+� ����=�V^�ޯy�E���H�D�k�+�=�t	Č�Qں�z+=�>b��@K:�Xt� �W�Y��,0qٺ*[y���X����:onº�l�Ty%�Ǳ��1�%�&Rg�+ ���1����B��Y�^��BA�v�K#�����N�`wש�2��*�[J(��
y" P?\)8��o�o]����%�5	P` �Ȧ����'0�+�dXw�<-]��m��:Ga�:/�/�O���9".p�h�S�OxI����>�G�d���׶�}5#sUge>����X2h&�%���E�W�N	7,ȕ����ɇ�B]w�gx�^ӻY�rD!>:~a�'�v m�/�.i/N�N�����l��h0��GIzj�CuZp��-)kJ�@�!x�T#/���Uu���Jb"�؜�}��Kt��n���#�� Ҵ��K��C�2!g�5��vJs(���L&x�?ڑ!K^�I��\G������Jؕ��2�5�b��`��\�M�qv�zb�՚!�9��.o�D�P�ft���D��H�Cj=^g(��<�a㒮��	wu��ĭ�l���}t	�6�%5o
3�3-�Tk�M�}����cLk̲��.���m���2�p���N��X3�L�b��g'�[#T�V֊�FH:4֍G�c�f��#�Oc��W����Zl��I�[N��ϞAvpf]\�u�@�L��9S~7}-LR'��^�	�����r�8����w��9�[�M�%�G!Ve		�O�Lэ�{3'�4�;&K��h��U}�4��H�vIO]�<��9��0�_AӕGx|��I��A4<'%)(2<�UŀR[K���8���ۿ�XO��Z�����R�^T�	�"5��h����}x�^ޭ�y�.�S�������٩zW�W	�Y�B|Z��|QP֍�T�\K�\����|ÍHnF���A��F�5��4JB0�y�L]���5"��"SIΨV�h*�s�{5�\�/�;��J2���U�Z�������W�B7��.8�!?��A~���<)5O+J����Q20ŵ���-������5��J��~���n�P'�|�p��q��y��.���P�t|(���?��4x6̄a^��WS��[�7��'&. LĞF���?���o6@Ζ<�2|ѡ5���뚻;1�":Q��'�]�h���!��j}dw�y���������ø{�KI7�in"��A"%�^��g��buCu,�c��;&-��=��r�}��n��x$��o#͠�BeW�iE���p7M��(yU�_���EIb�s���h��f��|��3I������]G\�g�a�̷��O��yk��=i5�|�z����5;LY�͔�x�d�-5x�� A
���)�V�LR�P�`{~���F<��.&1�*b"�TN����)��8�
�abL����=�p�)~��I4S
��L�x���?ͱ�U싳m���0�2�\�5 0-��\15��e_��+�[.B���e��ƈI&
��Zj��,�BBb�[�N��G%\G�:���t)܄�iIH�c7�5��D/[�`��y��S��7� E�j>
��ޡO�3�k���)�o�Cf�OH�� -���ܸ�L+��7�G��Öp�F�Zq�pti{�ɥ��}�)5�T�L�� �ua�`vp8]r?�c;n��=O��&��	%Ӄ�4u�1��li�g�bm�ss��H@�^`:>�0�����l+n><ϣ�����XQ��=�<%��Cq�m�5ּb3��`hs��� C�B��%�Ѕ`~}��Ϻ����yǗ�=\�B^��e
�Op��#%@��8f��$8��ࣚmf��2t��O���B7ȡ2�R�'Cb���Bcpא�=֑9:)��I��)��Y�"�E*	_����,�Q�jbʽ9�3l��$ϝ��Lc��-�1��~i�����u}���3 D�MSC�-�����Q�QyQ�� �ʄ���41��S�ᮬ��N!��SAm���g�cnZ��E#���9�<򝽕���Ad��<���f"&R�$����l�TYP��gB$��j�)�bɩT��c���SZ`�-��yRt�H�%�������b�X����lX�
�fY�w�_�*X�1��{�G���ɂ�v��1m�+�x��ˣ�E!�h����fM��i"�0%��瓠(�-'���={Gɏ��6��2�>l�s����a�ݝ�X�����쯜L�T��?�8j3��-4$�H��tFS�C]4
gF4�}�=dί2>rS]s .K�!:��ꄸ�=U�p~]C>gQŹ�SM[�n���$�[,³��a������ck��Ns�>�RH��6��+i8;fY�J�����3���w$7k�u�]�=�kց���!�׼�Vn�P���,@�7�
�A�ސ"�.�"e���CeU�b/i\2�_B��b{�ǔ��ʔ�y5���s�8��m�?f���9����,@�h4�5U���hҳ���w�p�0�"���t�s�*�L�AS��q��8�X �F�C�6?�h��M�3�xC,Z�	���^b(^q���ٽX�0���b��҂夝8�oC��;�(��7���|���4�E�
o8�Hk�e��1�5��_Ɉ�ͥ/�(w��'��D�����c)zʄ�lw�wZ��	�J����D�b��~ȁJ�Z�Q3L�NkV�P���@�_�{P0��^w�\�E�i}Λи+�q.}��/Mٶ��#8��y�r�nl[h[����3i_�֑�`}�1�;8�JJ$����J	�[�$c�O	�x�R�G��i��eQ�����h\x~�f-��:Xf����B��q�/z�D��F���ȋ�GX�����V��z��j��=K�&+r�#���w��F��z7L�-��9ѝ�J�P4�K���,]�uǫ �����[�s���d���l�����j�T�{�'�M�H>uR�F��xGЛ�;��}�T�YƯY���b��w-(���Q}]%b0! _>����vLM���6=♮���Iޅj�߼��V�����i0�E
v�̀o&�0���)������gl���\�483�tħ��[��j��r���?Zl�i�M�� �d�#Ƶ��f�����c�ϟO��Юy!sF�S�������h��$5c Fxq*��Ql����w�Eo �}���l��K���� י,wE�;����Q��_!���9��s�Eȏx���?2I��Nj��J�1���Y9^�
��'I�>�H��Q��u����E1�r�	ӷ5�F!�!g��6��a�d�D�cT��~����X��;��mJg��o�'5�?l��rN8.A���/dM{�e�J�&�yAc;���Iw��jG'w�S9�+��~�T�ƜFB2.�h��,m�3�.0�_���.W�S�?)�m� ?4p�]��顱}�=U���J\�T��Z���mg����j��%E�r�8�Pk�J?V�]O�H�� 0Va9���[|���Z�-���6�7e����o��K�-�r>�y����D�|����T��B��yj���8��������D��o�	̓�S�����گWU��&���C����-Yisb��.�f�2_�	�:
�N�__X@�b��`u��m�[}�m���l��1����G�;ti?K�t�4�!�xTar��EzY��י ����أ���.&���L%j�6�႟z)�$���m���X&[Ba�U�S�(<��M��-�ԗ���@h���C���h�0ԏ���aҍ��둒X���_�mQG��v;T|�E�� 0��$!�M���Y�])����A���8���8cx����I;q��­K�ȷsA����O��|��~X�-ԇ���]��֬�o�9�"�xT^�k\S>�����.��|OTp>�����IL��4mؚ]�"յ� \U05A�9&�p�~�?�e�glK7返rq���,th��՛б�4�Œo�'�<�*`����ƙ��vo�q������Rvic���4�c��[S�`� |������- ��$dE4��Cj����������X�甞�.I���F����S�zt�av��RJ��{?�uB���^g�q��������v6�&�U�)D��jJ��C��{@TF}�.��a�T|�lN�奼�t�3QӋu�T?r�/�S��� =yB�k$����v�����r+�k�����	1��[��Cn
\
,����I�ժ��Hs17��b��Y"{_'q���-����`p�30t���s4�Fy���{cf��g��_g3�6Y�߇$����5�fE�$k����� ּܻRИ1y{)�-��k���Һ�p�f}s�i�����%|��?�OA���8�I��r�����*^���UIn�o�WR����G>�̺4���~�ӆ���rqCg�P}���D��;��?�I	ap��U�h����"R�0����<�b�s���B�ήD�(��	����+f�'��'w�˓��h8D�0
�e�%����LM���P$	�^���]���}=�C��w���1�F��V�fTY���c���x�ħ��#���S����q�&��c��[gV������ƑR�4뙾�m���?���i������W�7��x��W��#�f,ǭ�jmL���̰�T���zߋ��'uG�KȄ�;y�2�?�P�'[�1��Z0{���=�~`!�_jb�!Њ�j�{�3�:Y�.�d^s�U��C����-��c��79X�����N���m5���8E�3$�bպAD�h{e���
	�ܻHv���ӛl���>�#_/!��{'lgS5�B�p0�a6��^�N�SOEw�;b�y}��I�� �`�;/��rˉy����lp� �N�����IVq�/#�\+�|l���gZ�jk��n�ZC�t "M��^`4f�2_�FY]����~�Uw^"pܯ��f1V�)W�L��0����[&��Ҩm��f������3��U�����[��d	*��q��VMc�8��
�kĳK��1N��i��)ߠ�����	 �%�˦@�4�Sm�����n���L����ݝz�9�Wyek_��(�:�$����wF��b��b�3!��QmFk�,�ZyI�>	&����ȼ�F���C:*h�,k<�4^P���g#L~�t]�~}�ĕ�#$���i߉�H�?�k/���F���x�n'E�#�T��JKy�T�U�p�X1]p|���_\W�^?��x���:ѤT�g�w�^c����yE)��C���C`�o����|�Ni~��K6&��=2ZN��k%��\�|/o����!�W�r3겻*2�"������z�D+aa�����ܳ�w�e��m�d���̘�[�}:�4+PJ��K�76L��Rp:`*�X>�p������~D��sH����������V0��Ls/<�w�M��&���a�Jy��栽��� &�T�"�@�sƖ� p~���%[�㺙��H��ϫ괹��+<�J4�B��.�J�e�}�n?3��@d,e,�e�4�.I�����u 0nc����c%��ϧ#<.��L�%
��+d ˲m-��]�+L����X��M9eiĠh�#���=����X��Ǽ���c�w'#q.O��h������0e����d0�e0���ΥW�ç���f�F�B�KԂ�e�R�c׳��{Z��|ߦgP�މ�
`מVTg/�M���t��y��������T�/�]�X��ؿ
�U���5]����#ρ&"L~"x����2�@�Y��h%��2�s)bN��~:���>��}�R9�)Ue� �~��J��V�y�AC��x�u�"�b#׌{�����l7x�^|�ǵ�k�|��,�Kc% �	��?����Х��̽�JS0�̑EG�&R�����-����3a0����DU՗ø�Nb������)��0��� �����Z�x��2��Q20�X�2;�ꨊ�o������n|��i[�]Ll�oh|^# $�ʈxk�ޡW-B�#�+Ba���A������u�����]��;��U�_���eq��gF﷧�}�Km���Xn`�;����c�)�p~������U3��q��f����]Jg����M�v�K+��Z��e�n�S����s%�I0=��i�m��� C�
~;)w��*��ĹH��
�����a�|Es������
�9��b���!���O�3x��q�[�|4��Z4W����m���Ưb�~������3�W7h^�D��M����6	�U�0Oq��%���a#	��,�Bgj��Q��o���XԀ8�[qOr[P�g���R�#��̝���6� �q�Wy�UuV�v�,WV�����N��Aq�\���'���f�����6�?
𵭳B�Ԝ*����˽�ݎ���V���=&dH����������,Ϋ4�����TV�o�����8�����O���s������S�z���-r�>�1,4���/~��<q~�^Bq��Y�E��^H�>���@�ͱ���J������*a�X��)n�DN�1ʡDO��8�ێt�n�-!�{����O�n�B�-i���ǁ��(�W�	��b���)35X^:��Fji�2�p���".�(�]��WR�k�8�4����=IW�E��0���|1x�bD�no^�Uj�Z��m��/�)�R���F���?���ZG�E�����N=��3���z�L�"j�#��!W�{\��]����9ޭ��f���B|�_^��yRmd0C@�x�3���Л��2y�wS�]w����/XI] }���ɼ�>!�;�"��73"��2��w�@}{����×��H��͠{��3�뚰�W�f���9�y����/����6�L@�\^�z�S�������tm|\���x�,k}
�.ۗ3蹬�6"	y������Ύ� ���ĝ����0y'�?s�x*���̯'P�a�#�,w��
Q���5��ro��hC��?gV���O�
^i�
~��*�:�K��Iu��M\���;�,=���f�a_ʫխJ�Zq��	۝��2�:z��s�eT�T?';�&�IoC����J������mF�eAf@�孺6/�o*����k�����6�(��2�@2�;�ٸ�0����{�B�3�j���v�q�R�X�o"�+Ų�#��W�̆�X�JE[���T߶H^��CX���h�=�j�a��P;��� m�c��K�0W�c�-l�76�-�9��� ��������G�����&`�3G_�V��?����do�캱�S�D^�]j�Q��z/l���5E��k�Ȫ��=U.�%�뛻��g���+]6���|��)�RUj�lm�_�..���t������	t�;~p�b=:.e\qժ{W�#�q1�eN�<�ǁI�Ϫ_c����PGOp���?��'�VLZ	�V�ޯ���:{]�I*�d����u���`��3o���r�T��1��M[6%kuQi92�o;��۹EN����a?��}&��bx���@����er����۰^�]�ˎ~(�K{��R�S�*n�fVO�Sa
�]���s�h&��XG8*��ƃ�6�M'�+���"q����H���VP21�s޿2%_�q�C���`6��m���5@a���!䴆��SB�-L��gM֛�8hV?��;��2*L���w�&9r�w��xL��q�
b� ��A���>FѰ:��2?Bo��$#V��5$�>D5V���C�kМ>���z���#8baB�d��8;�-\�jE(lW/ t?��*y��D�[b��s��2UB���O�ט�v�����l��=ܺld:CȦkf���ˌKٹg�@ǈ�@�6g_�7���G�Y7�@�e;�P�RA���z�vI�l,.6B�S�����y�V����B�����9vx�4=1��1�Jr�tOT�{C�!�M62�y�ZeW�_�;�k��.w��:fӝ�<ߜR�:l�n�4�E�~�H:�@eM &�"ߓ��"A�O�_����㪔��Z���dޔ<���hlw|��+��na@�ݾVPR@�j�9h��ުZ������p�4v�STbp����l�t-G���x���ޓ ����wm/��9G,h6W�& M���;oz�[�80�iDHp+�����(��W�۸q{=���� ���,�|��=�9���v�����}������\�2`تhc>���H��Vx}���6���*58Q4��ɪ�3/x�Q��l|�o�ݍIW�O=c�xs�|@�0-����jj����S�W����Y�~.l�{&6Y�y���T�N��n�̞	�z�H����=��u,�C-�k��>J ��?->��Z>

{^b�S;��sN���Y��D�69
C?2�t���猣*y]��}(��Y֪���"V?��w>^r�Q�+�Z��i�
��<5���~e2j	��ʒ�G��T��`�F����r�5��"op\@Y�"�*��ǅ�o3��k\}�xp�aO�܃Ъ���K0����2�, �
W7:�\���f'G�Ċ��$��a{l_"ZȵG�ъu�� `�E�#V�Y;4uY?�~	�`\��"�;e����;�Kz�P�Ca@#����?���j*����g��)F�J���|��@O��v�l O1:Ğf�7��Q�;ey��x͠����=i���]5D'J-�F?a�78j��lvO� �8���9��Y�1��|���D��R���LbH�rk�aǿ#T�w��$��d�\�pcL��{�1{�FW�Nˡ�2� 2}�h6�9����]�����8�-����/6���&���Y����}�[�c��]�\�Κ|0�Ҍ�@�0(KF��m�q���r¼��,9Q�7�A��`�D�\F���6�)�Kiop&fG6r0	w
��J�5[�1&W̱�Ho�6��71f>,����+�޺jI�H�S�Rvs�X�1��E��"
<�)�h����~����v�Rk0Rz�@`Yk��Rw�5�(R����`������9�o � ��éU����%tSL�	밠�h�;' Teω�ԯ�8�Uӝ7��u.�=��>v�����>���}�%T&S��s�$�1�νE�9��M>����Z��H���N�h>$=�tj�~\�+�(�!�J��B09+k-�n�����S!y��~��#�@����[H���w�\*�?=[�����﯐j6~�Y{ᶿJ��R��P����'K2*pH��	����7��k�\޹�`�e��TQX>�X�/qX�8�"-0�6��_� w��̺����������Z��\��q㓓H[���~��P{PxB�n���^D*v�pN��.��{�X|�HP����9h���q�9�;ʂq̄3���uU�r0��s��2��ս�u���/�o N�K�2az�����ǐe���o�ǿ|J�unM/���Ȓ�"O�8�+`�ʛ��bUr6sĦ�\'��9	,t��2#�L�$G��2ģ7���Χ�&��>G�ƠR�����+�U�)
���ҚiRv�Y�]��O�f�i�`�����e�1|�3˽M��嚮��x=�R���SW�tĴ��%_�:��;���e��ͼ��~�<¬����%×m�¦7K{���:qj�����h�ȯ���	�5��D`�|)�T�,` ��u�yU�G�ì!�1�&�6��?�]�[�0`��~��o�B��r�J��Ʊ�-:F����cOO}͇��?�	O34�w�p���dB�������k��ӛ2+h�(IU|C{�>nb
o3%oD��]̾��Ƅ��Լ��
w����ջ��f�@��Mb�7�k$N]��C�1�9������ (��o[PCN-��\�`�1��S*M���:�ݤ�4��f���$'�Ii�>׌�^]ER���#�?�5и�̲K��z��*�0�?Ã�
�+�'�9@�'��'�է)1�ŏ��v�/���B�(���8^����L0S�P��f�?':��I��i��\����L�Hz��Q����4<�c�������2�c�N��9T��>�Lʬ	�� �����B|��H.�OUb��K��/ 4����K*-�Z5��oSĤ%@2����{DC&(!2.&��z�2~�i�J�0�X���k7�ؐL��M��o³MU��0Q��7y,괈6����Z�#Ë����\`�%��o�k
!h���F��i姭j�'�|�'CG]���P��>A�f��������s�͙�T]b6v�t$n���%����.���lr׍&;b~��Ω�%޻�\H~�����jZ��K�w�p��v0�<>��/P�{��M{ �_����:s,����OJ5ԗ���4���΅U4ܺV�:�g�W\���K�͹k�w��$zw��
����~�+���"�pF��4��R��EY�，�{���zp1�ނ,p�F�t.b��Ke����BA]m;�2T�Of￶�Α3m���\��E��CR䦎�d�C"&b����O�M�s�3��߷�u���`}��}I7����f��?Wʍ�v�P��w��T�z�g֦h��^�t�b����c����
��T�D�����/�*��4��`����ұ-� ��M�5�-/zĚ��?���Y��W��O*gQ�3�y1�J욎��/T���ȆlApV�p�v�5N	��ki���s��9�����h�^��]�+��//�<׀���+����(��Q8k�O(��1�Bw$p����e��
s9k^/*�ċq��Aa��]��$g�0t���cp����X\�+����pV���9p6d�	�W�G-�[ W���lBv�x6_�u��հe����-it�v���Q��Wj�@���ǘxe��%)�(���>L�m!N����p�*p��L�W��l�U�r ��9�6��}�D��Z�7��]���7�&{�J����q~�>�;��@�`<踯v�anV�|��	"1�ޡ�X箜������_����!,9���oͺ��_e����篟Hvc�|�[˓�ﵔޞ�����-9�Dn�H\�Am�Q`�ȫ���L�ۃ�6��Q��涯+�(yJ`D���>�j["D@��O�#Yמ�*�7!�b�F�=�F�$_͒��~qo��@��0�3Y�������:��������8���#ES�����D���&�G˴�c���1�\:�����u�R�@����tz�U���u�m?�����#߄�`�U��k�^툏�0�Zl󑁸����D��v׏��"��Bh7k���1�-���8<�e� �YJ4E�zn����q��@J�-�X�Z��!z���v[���1{N����yr�s�!����H���ڷc� ߴ�iB�ي����p�)�Hb���si��aZj�Ml�.�G���H9����z}�)���� ����fW{�v#�����=@�i�W��dX���f�r %���3v�Gi$����)dE+҂:�L���-<�/�WU��~9�p��Px���Le`:��Vn�*�BZ9��v�'� ��0U����D�H�`�h$�_�p��W��9����M�����h��i�(�ƌ6S��䨚���$�]~i^V6:p���Y�A���ď��[͖8��|k�}G�Y	gV��yΏ�CNq���5U��eLs��A������ƚd#����'v����Ie'u��L\���׍V a�m���/L�(��Lk�v�c?�H�M�H*��k&�D�c�}r��0w������Qes�w)1A­^8lsV��V()g�8s�J&ݿ����濫�B_��p�V�T'�"���]q���0,0*����=	m�W�/҈��U8̎���y�b�p%��ґwש�E�Ȇ+��_����Q"K?%��Nk�����8�68dz�61~�T�%&fA�C��7�5u؉�~��lY,��;�lq����WI���"W�@4�U�bvJ�~R%�5���j-���-��y6��Zܵ�}�7�q���WJ����GI���?B8%9p�*�0a1aH
8�y���T�Vg�<x��8z-��ph\�)�_�й(����(s�8"͖�=G��]����&�2�VUZ`nK��J����o��(>ťI@U�Á�=J u-�Y��g�ǫ�tkZۜa�˹�ű��]��
Ws�1�0�̵���ͬ����}
QfQ�s<�ݭQҮ���Kq6f�R� �h���Ŋ�pu��9�����*�R�|pvh����3�|q�]@Ng���i�K#)e�?4��s�������]p�Q:v����%J�{��������� .���o�D��qpS�x�Z>ʹ'��a�JB�����
���L�^A�č�2��Qy�!p��j&y�?�ǋ����+��њ;!2yZ�>�40=�M��֎�/�t�Ey�w����k�:�Ί�d�1���F��t������K�k�ړ�0[�ʭ����v{�>@w ����UX)%��j�Z���Oh8M\<b����յF3�)6�7b��ړ�wWlh<	�ɵ���)�T6y��fW�0��O1�c��O�T���H�$��j��`e���cX0�C]g��̩������)�#v���x���i��3Z���T����h^�-{����E��q(��IB
h����K�"�� ���f@G��{�[6.ڡU��DF��=��;��ڶxe��p�O���,�̴W�抵J^GQ#�P��U�=�oL#)�FR�D�2RJ#���D�%��������<�����K[�k���P��-���q�F�Qk۱h��8'���x6�)������ڣ!���x�j��ԋWs�Z������f.h?�Y�@�Ýx�0�Y��t��g)��ã`uS���l]�i"�&v�%P�.6>�c�� ���d5"�Knjڡ��S��T�݌��Ѵb�A����{�m̑�l>�`�ۤܵ@�H�Z����i98��P���չ���ԁ��aw�����z	YCE�����j���n��`ӛ����Uɂ�gnPk�����S��`� >:�r	�;�Ԩk��Fڻ��J�����g@亮�1�ژլs�MH�-JVc�����4��?�~'X/��k�z8������	0����_��,��e�V\;ȯ�+^ �c�R�̄��$�?+q}�H;9\B��u�*�����}��8q��4��gH�f�-��q����\%a�xņ6�Ǿ\kɼ��'�B ܀ئ��b�a��^�X�9�U��h�ፋ5;`�P�*�a�[T�����>�H�r�Lm���]㩍�E�>�F���`�C��o��� ��pa`h�_6�6�r/Ll���dv�tE���9��\��2m$}=��咯˒s|�,C���
�'���ʍ���:�ٕ B�Ǜcf��H�^�ꡆ�	�\ gڹw���ݠ��+!a�AL��y�	(W�Vdm4��Q�r�(�i���6D0�6Z�؎���J�j��qb��ɕ��:��݌���s� ��t	�^����؎�+i�凑�$n����dmQ!e�vk�jl�'��'Ƈ��M~hO�T���p�F�k����ᬰ�M������o��&��Z��7�]����mʪ� �u�l.�N�2�ߢ4&��1�]���!U�Tb�JY�~P�X,�lj����?����l~�}\������(��pNTw?D,*h�v[8�lI���-ȡ�&v?[��y�g��|�s���7>��
;�8�"0Y�TΙ} �,�TGMe��ک�FQ��C��sm�ZyN�g���
�
�`-ٓ�@�?����7N}˟\�aA�659:�������b���/�����paU�����#q��`�E��df�>�5���C�н��c��!S��p���A��ǋ'�E$������w.��2�?@�`�����������C��0�i�w1?��� �3���7$�
�\�xKҋ�+Ez)���ݖ� d7����4`�"Bh/��q�1�`h���4���>ʥ�S}Ź,{�Jau�߇�S�f�r���~�"TF����/oc�p�ink�#ɋ��b#觫�XfI�7�ƺ"�}��c�<������j�k^���� �����Ur�O���JCa��y���b�!��)����]L̋��]-�.f?�U��u�;
:h\e�@YP}����)|�=�y!z��Za�����e�xWJ��I@��g�>$'7���Q�4Sv�	���C9R�?������c�����2]5XIδ�T*\?+oE' ��������$e��nu��7�c��cg�eD@���P�B���!�^`��$)oo_��P�L�,PG�R��M�F� G�k>�F���|���L�'��"^�.��M���.�{p�xY���������������ĉ�f����^t^�_V��!{l��4�ߍ��떜ܲ4m�TȤ�@�����̩x�@l�\''1<J7I�o�r9���鞭���R��?��To9��ֆ�@���Н�9�}tD� EI�{1[8R�,�˄fv�M�,kQ8��+]u_��ئќ�Z�Ԃn��OAMz��`����1��Z lz_Qt�R���&�z���	�?v�� �f�?p �|P/�A���0$����"����:�	�A��
P�-����+w�-�(��}X���Z�+-E�U���en�2~�O��fo��z���BD~�77Y�Ԃ�F/��mު���i�����.�6AG�����]��F�om�k@wmq�贠7�8�DG�]r���\I�w����Uj�0�3���Չ��L�iD5����ৢB��%�ظ�m����jf��g�ʐ:��yc���$D���'#�kPA��@J6�Y f���߮�_�;����J��xv��Rwk#>T�༛
nqs����b�$��琙?%�x�sؿ�r��H|>��2�:�=�g2,-��-HJe���Q5M��fA�=��>����QՓ�i���4���P�ٝ���������0�6��c-�������s2�ݬ/Q�l�2�=Z�p�`Z)�H�)c���F��n��Xȁ�����(�nZa�O�F����FC2��eq�Ax29`����w�u{��N��`A�k<�[v@����>��t=�I#fm�D�.�U�F�[km�v��;fWi,�)+T���f�����b�.���tSH�>�P� gQ�,§h�#-�:m�8�.Ĭ����b���p��f�Gv!lӮ ;PE ��P��0�A� ���sW��<��b(���"��Y꾃։0?���"�`��+���[��U`�P�ۘx�/X*��M7 hRc�?~����_\��ETr�v�#��2�Q���i��
�]VXE�D(v�'oC(rd�����Z���t���KcG's�^����%;!�N�R��Q��d!:�i`nm�g���|�[�K�r�<�hb�v��{}QnI.��`h]���I��\��X6�	�\涴�C7��[3a��S�$�	H-T��u�ҭ�����a�MSd��}�B��!�C<ړ�T��I�<o9@�ο/��=ǒ��2�^��RА�j�����X3��}��/�?ߪx�N껑wc�&b��R�����,��J��3۬���ƍ��yDq�}"��<�ܦ5�Xkps<V�"�4j4�F��������*����/{�dB9�Ԭ�~���y��b�}��E�%��;[�
�#�"�#Y�9#�Kܕ�^J�t\��Ɗ��
���^�
):G �.�2�^���qJ0������`
�fW�}�;ݏ���uZ�i��J�Ġ[�y:2-=�	��'�U���ё�L�C�̔�n����G��SQ�:D��C��Q H� ���xL���aAU�r�l� �(��p�7t]�D�K�a�-:DD�{���=z�ۉ�a���uF��׵�0��It�Z%�NL�@3irP�;&�����\~K�{da���lRt[/�d<D��O�,��`bB��¿�YZ&ڠ3h���>�΁���g��m�n��UN�qæ�`:�ra�b8��$j�P\2�� Q+��ۄ�V��Lt��f¡1���������P�R�ǲ�g�#�6q�ɛ.1a�w9�ZaE�n�l]�pO$�:���6�q�`�Y�е����\%:5�'J ��ؚb]m<(\>f�i'�R�'&�Kz�o��M�����Q����
�Cu�x����a��x�|޿�b��?}T�1�Y�?�!�}�7nV[u'M�IF��z�Z��"zh��ly���j��%�������V�8Y��g��9�!��~�N��g��!�n����j��*�R���{[�&�|�;�`Hq�i�|7Ʉ"�L�����g���x��t7Qq~����>Y��-)B��K���;��[M��w�E��8ɕ��Y�����{q��ɺJ9s=�.,@��tz���$c�Y~�⾵��K�r�r]����V7Zh���"��$�þ��z�C(����<��XN*���<�����w�X;��Uɧ�� $R�����=��!p˹��Fg��¡���9��]瀽�E����&QV� ���r�(+,]� �E�������_D��T3c�~�y���������%��i�|r������a����h�d��p�$;�W2[�� 7Dg��g�����^_}�{�0�"���B�w�$b��bY&���nZ����{�i��3^u%*e!Ox���ا��ʐ��n�����.�BGEŭ<=�Z��A����Wn58\�X����Α�7�?:ϓS`KN���Wg�X���+�/E1���V��i�����rS�D-�>4d����i�Pں�+@��Ƀ*l�F��l~DFI�W�����qb�^v^�X|8��B畩j|��6�QCRi>�r��hgr�z��'���3���~N�����Q��)$�H�m���t��H�3+ߦ���y��m��?a��f����)��0u+;�F>Uù���ʠZq"m~a�O�f�a�n�]���*��T���Gab 6�'�_�7/}���{���ፈf\#� %�������0�p8���s�%Z�[�D��- ׬���-�'	`	�t���9��i3>B���T�Z����Y_���Q�o��^KV���]�yL�L����)��>{�ۘnJnf9h��J��+��gנ��<#a w���ȅFƯ���vA�2�]�^��޶?9�ݎ21��)� O�"
Z���D�����֐�¶ـ�g�%;}��
B�5�Q�+�q�6"{�RZ�;�.>�8�R�2L�v��8��HI�a���q����۷���d��P�l�c��Xx��A��z�S����L҃�aj�)6IH~����\���W�:�YI��C2���1I=���T@)�M��:B�O�j+�����"�]��D�x�����B�j`��|��l�{�a
ȧKh�S+��	O�
Z�ߜ0�Ǉ�_�[�a0���W5[��츶/6rT %U^�lz�B?^���[���P�o�襔�MC즭�50��ȳ��)7@�-<lB�N�Mݖ#��v����`�  �p������^M/oL?d,W��Fٗ�ϗ�j��ް���Uy�)�������Lf�Ќu� �;��H���l^���k��<Kt��7�
��@�f&��^7�A�
�'��X�0Ax[ZJ�;��cqS��Vʙ���\a��1Z�qkg���|�/��8��ۄ~�W����j+v�+�{���5��ْ	X�Lڬ�Հ|*Z�!��m��w:;
D�m����4G"0����S��[�@��.vϵ,7�鋚��i�o>O&��1V���O�~��F��Y֏��kIᜋ��-q��[��s��� fYi$�zX��I��6�N[`�)�0���^Gb�8:a@Ϟƭ�7d� ={���$E}e{h����� <]����z��[�V��d{�H��<�!�!Ħ7V�d?���p������|��R-4n���I�-z�=�^B5R4e)<Ń� �|�4��)�Þ�����_ّ~�!F���®o��PD��G��;<BA������i<a�X�oVf��~p��G�������r�q)˩�1�����Q'-�Hw��\#�xbsNaAN�Z�U",�#/�%�~�9��<���Tr���(|��,�K&�?s4�������0Z�S�����Bs@�&�(?������x�W�wY�H3�}��N-������.������Mӻ qZ���6����~#a2~��g�"�T���IF�0tH'����E���H�7<�����������t�1V�Z�"1�<�Y����.�C�z���o�X8;	�͝
쟕��餭h�x�i0���F^��9%���ߚ��<��9�%�=��v	����:��s��u��	c5o.b��E�?J�1f��t|nw��J7��(0��'�N�XDl�rkd�H6W2�6�i�{Q��,z1��<�ͅ��Z�.��,v�T��E#�i_��Y=U�ou���/�s,�Ѿe:Gv�X1����!.j��5�#5���D�e�#��M�1����T|/:���g�3Y���K[��y�JG��4����9��������29��BP�:X|C	h>w�Q�r
����F(�?�C���U�߁ݮ�Ǵ� ���%<����NK�cߏGRu�@:�ғ25�NmG�Ʈ��=c?���?c�����wނ���������!�������O�S�n^I��'�h�q�6�Ü�42����"��x{������Ա��	`e���)�������<�Q��n����U4o�I�Ay7u:E��q��Н�|].���QӁ���,�I���Lޯl��ة�0��)>��tJ\���@xS:�q�i�]���:;��$;�6~��ƻv�e7���U���g~�LXA͜T�%��J��`&�1;�ˊx���5��]}/'���}rZz�NvY�I�?!���TxgG\�����������eװ+B�k3����Z�a �^��3y����M�:�Ń��E�e�5��Q(m[{�az�l��N��N)��J�
�Ҋ�^Ԗ��&��a^W�����FfB]�h���~�V�����@���&�m�v+l(,\�� �h�������E���V��U�QN�y�ШL��Sfn'D�y;G%�w�4A�_�@�Mڿq��Fhul�ω"���ʔ��8~~�4<͕(j��'�א ͰI�,�G�[̭H��������╛��-g1ڇ�p�f��m�+�#f�?���PH0�,x�e��MD�� ���(������uMs!Pm2��/@8F�����N,�?i�`��6�xZʋ>���j�[�_�̺z8 m�C,  �e�fLs=�������-�?���������9��0�z�h#��C�v.�Qb�k�F���� � ���}X|�%d��߆T��Z<��Ʃ�ƟN<rC��B�û��A�5+�sˣK�#ь�	�)�E�Da怐�f�6��_{˭UI|�a�*S�|I2�9F
�r�����MVe[��#e�Td�Q �ll��Lv��������EzBj��#H�R#��L1���]k�7zz+�}�N��"a(OE��CcRί���B|w��٧��j1�暉���"R�9#L u	a7�`��erD��i�-��Я�(���q������Ǌ%��U��4�z6	h�p��e��&���:aw�����Z{�'��6��~����&��/�w8 \�$*�+k�W�d
�3�-��Ki]G�M~�h��9�G��߼$�p�ϧ�ބV�?��D�2QA�3�^J�'��UN"���o��KE�˞��+���+O���s��S�.���A	�\�����cY��&�3�*B��M�_C�X�=5�Մ�����*;�u����/��xr�҂���#秩	��Oa��?۷� ߍ 0��Ykd$Up<H�E�#�|0���d�ԭ�t���w)��^�Ji{��Ԋ�А���3�5:uC=�<�SLaӆ������i�	݅M�_+_�����P�fT(ƍd�E�` u�?˼�o%���b��T��u��hc[�=e�:�R1۔�Ղ&�t�	��q���jL|� �qY��*����~���TIZ�vdB���� ����Wa�����es�%��̩�Ź	LZk�d����^�"����&&��8�\�'jg���q��t<�e?{�ӕ�|��j�?E�D��~�&0�?���
��`[o�%K&�XhBM�`d��ʥ]@��t�&�W�#�B�0NfHh��?v S)%P�~&� V��ѥƤ�^����H.r@F���_x����F��>|�$J7�)�����Q�V��$��פ�Nw�d��T03��&���ǘ���K�fKڇ�#����ʗ���xK���F���=�UHT�s���|���$Ll���&�<�^�m��J��g�=�eX	�?���-�޳���2�&*�8t5��d��-RhZ���zA��)�l,��/D�@��}�����Z^S�R:�^�ڝ
�!��ppp�>���xW� ʛN����xj�H�~��X�&fҕ�C�|�!�/�bD�[�%F���)ӻ�n%����oH���8Dt�N����~Ҡ�T�A�* 8gpͫh�j
�sۡ����:�ko𲝆_��=�\l- �c�Z�O�BW����hJ�����&��W �o��>r��[��(��!.��� ��@���3��`L�q�JF3�R-�a��ܡL�p^���傗��0�����aF�H�<�6��Oıd@�F|�w
L�T�h4�)> �o1E�9ߵf�*����tgK�)�?�w�� ��<r��IÿK+B���W�b�p�F���c��4�����<L?������.�|&R_�$9�_-N��c�!Ay9"\�ֹ��f���GT_̗�jrPS��$)�Θ[��o�l�H N�Z\�B�q���q�ƀ���C�T1%-�4��G�T
u�ou�]�Y�[`q[�l3��ԕ5-�'�����Y���@����}dbM%�C.�B��VF��p�3`����M\,����ykc���Z����+2��E�vEl?�ҌU��=�,˞d������;�*��]��:M�E��}^�M���>p����+G���;<�:I.�@Hgb�UO���Ma@���Z��t��o�F�ˊ�V'�0��!�F{���.>&�3kt���n#��k��/�U�/h%BO�y����| �ND��Ԑ�i	�t�J$sz�\���QHY������!:B=�p�S{��"}���zz9��k�Dj�������F��1�Ӛ��^J�C���?��@3�/M�QqS"�ł@�sN�`��"�Е�{�|�龶~����n��&��R�j���HU��qrAD���b��b���z� #ɂJ0�r�3r�r�⦓�h�\'��t��H�z�Dwm�O��	��yt�Uu;4��I�{�������D%��Q=�֡�z$p��=�:�|���Ĉy�S��v�3~K0зRu��_��H�qb��b���:�N��g�'@7#�s�h��/�s���=6�9�L}���:C��G�j�-ot(�W�/��a�w~r��WF]�L���sXiob�9c�Xo%�U0WήU�%��b>Q��ء��:'�eԦ��KY2���H�(}=��)��ŎK_��@�$bi�����S�q�h���X׭RDm*g$���(�,V$qƘ���0�X�l)3.�/��G�D�ͪ�
��B��ZA,
��UExa�aΫ��}��<�}T ڕ�i�h�<l&r ������ia�P&D���=$a�FkC��P��x�e�p����ͅ!�N5����Xj���x7��@�4���3��G[<�d�����;Q �����$�L��a:Ļ�Q����@\��jو�^j�g�P�L�f���\�ax
�4����8x�I�FP�a��a�!��U�3:AC� �5�|�p+p��x���@�uaJ���M�	3��tŞ��J:�Z�+��f�Nz1%�<t�|l�DV�����:��r�C \��=�&��4�� rA[�1D鎌P�'Y�)�����sȋv����q�(*�4x�Z��.'a�/�`3xBI٩�7���nK�yæ��������p�
�۽����#�K�I�\2�5/b
�y�]��<D{�z4l}ıd.��S�i+�~lHq>~�j�֩йt��<���l|,k��8���������D�I����A�A��<t,�=֋�S��2A�����2U��8x^�;���	�W�;�HJ���4,��6۰i����4.����ϟ�K*�b�%+����bΘ���j�ٿ|�ѤH�19:�tn��p�A�h�,�Ԫ�n�4��U4�l�А��A��EĨV����e&�ȅR�x;7���,=0ظ�t���-�O��x��{�{ zY�\p�\1:��"�I�c���x*NSG:fU�����bK�s`�Fl�[�J:�c�̏"����8E1W�	�v��i �<5?e�+Y�D����ѽ�8� 02$���X}4,U�v?����
�j�,�.�ho0���L~�����o���������󔸡�q�>@�A�^ �aOIU��AQ�`�ƯT;�n�v�t}�HV&�ϋ�}�������-Qޕ���X�l׺r]�7{eչ2���(��#����i��-XT�IX�.0;��h~6W�{�p�)�m�Ub���Z�4�>RB��!�Pm�~�o�	H�,��1�?����C�kb��j[�?БI��]z���l#�s���Ze�S��2�ls#��Y&��c=(�1�l_ow�ee�'���t�5�@��Y�P��Z�pN�	O5��UEdl����$o�K�g��gQ#4U�1��%��Tn,��G�;:����Z^r�G���9�DB���?0|r�Cj��R�놇-z�H�-�T��:95ķ���@��6�qBg�\�D�s2�̻@yO��R��-�7���Ka�&�n4�CD� ;8 >�yrw�kl)H�F�̆1�w�q��*-�ē�ú.��WK�W��X�R#P�(B���J��ӥ�q��8v���e8���DZ���P��� ��s��[�RD�{��|c����F<�/�	�@52���1v ��I�C��ZVk��B�p�N�t���+Ҧ��Mqh�VF��/�"	�H�f�j�����5Z��hcW�ㄷ�`��R��iXOz�v/"�!��}�̧�W��$�[/�h���n�J�*��<�l�T1�r 8 ��,+U#S�Hc���������{�HN�Cq�I���e23��Wౠ	�JC����)�6��FB��>�{�w-���x������4����CXg�yr0�v|;Ğ5X�&c�r-+ց�}�'�ȇ�`��.2!�iW��''`�M��Ґ^�8/9iC��\�=�ʓ�NɍSN��Ax4��l��R���MŜD��S���@%z�{�U�H+d]�"m��Z�C��:���I#� �Ϊ��I��~-����Bx��[W��έ	�4T�3�������#Ӝ	��O������t$��.,u��Y�K%��hZކpWx_�T�1{�vt
�w���6qKO�~ ��@���+�!s�6>�ʂ�_&$�RY�����y�V9[�%�#3_f��̓/@|J�.Mo;�%h:*ײ��G?��Q"�DϮ��u5��7��RO�劅�Hl��6��pf���Ӄ��s̨a�����{�Mc�.^���@�qP�=�M���f�*�~���A��+K���x��gJ�oS� �Yb!�qT����r:�;�!�;��ux�7D��,�}	FdXl����C�{"��x񇢱U�]���g[&�����H�gX��,�>q;��J��Λi�\���G�^qZu��7�x¡�Vվ�0�7�?m�Nū�
^�:X8př�$��47��
Ѕ�x�W$��Ƞ�U�*��GE|H{��/&v�?�	�gCɏz;5�O�$��}�`�5ܺrܱ�DR@�ᓻ��I69���I���x����J����Z��v���3!��P����m�����ֵy��� �/-�������Gţ���OL���̖�!��GjWv2+��hM���H"�B���]��aN|2�FD� EV�s;�S�n�7tƧ����������6iSu�5�mҜ�`�j��\A��6�*��0O?��;q¦��/&�ov�V�rdj�w�X�Uܭ4�;,��+�y*�������,I�!���i���O>���~�24��V��B3ޛË1R�������C��	��<��[�r+kU�u�����C�y���Ռ�zh�@�6��=�3����K ˿Vc����ӉNI翩�'AAHfcr#�٘�5���vZi�	�}�9CY��o���K1FqԳP}V�}��l��M^%�H�Vqh��V�1Z��*Dj��Q	�ƃ��*p:���m���rIkk!�`5�����۫솪���"�$��<�%�
�_0��y���{)�)[�C5G������݃���7\ P+#�����~�����N4��}]h�+[iv�q��U��'��_
��	���͸�I�>^xڇ�3�K�F��[����ӐC��D�L(�['�8��I���GGm���!�.�����D����ݐ�>3� �	|KZ^�#B�����x<�ٟm��}��� o��PG�f��y�t�!�gK�ѯ��K��v���2�|K��:�<K&��V�m��)t%�)����Ҙ;�$���%�4�3��k��=�������fJ=#�K��f6Ϳն׳D��T�ޮC��k���md/}Ᵹ�7�N�c2���%q[9H]�c{kC>Fk*O�""c!6 ������Ơ��>̿�s �<��W	4�~�7�GV�����2��&*}�&��~�ޏC3w`Y���C~��%/�m��}�d���+���^Xh�q�Z
�S�6�k�䐅��j�N��):��ϘvyU ������I���=V�U�)��t���X��h����1�% so�F���!rC7Iʶ渗d���Y��}*V���|��.���'�0� ����d�2O]�q}B6�]�Ѩ���95H��pL�~҂mK~tV@���Ɗ��j |GꐀbV�J��W��D�$�r��}d5�����cR_��p��Ŗc��!���N�`L�f|�e�hY�Ԫ� �ś�8�(�U���蟊�_eI�c=���g�$���ǫ��t\��������Q�V�U_�-{[���¾�FTAG�0O��Fn^+��ͩn�@]	��8�5�G�
+Ģ{@��zB͡��,���\]�ܤ�=�����B�pW��,����u#�T�*G*1Y3������3D�HJ&;���v�!�u�A)��6�Y<F�OB�DIl��^2��=��+�xZ6�6sc�O�սί~<ǡ�����e�1R���H���h�o�����nZE��(�:��-�	΂�g���2�X�Q�����苽�/ȳ�7W+A¾��z}�ϫ]�R�>Hbva�t$�5��S��?`�0�;��t����$� ��S�q1A�,�� ��%���7��������GD�-B����֭�U�����r��,Z
�-�ZX�W�N��a�"����^")��?����:v�(Q��T�-���J]x;�UV�	N�z�r2��)�L�e;�]��%���9�F�9?��l\���|+�����r�����ĂN@2#xD}�A�%��;γԞ�bA=��7%�T6�
���'Nu,[wGW�n^IɴX��	ƬN�k2#2�֋����W%N�L�I��6rY6p:�fq��������2�@-A�1�y�
֞��t��&��qCkpTC�~��Fަǧ^��݂��{bZVspc���#sY� E����H��t�fĘY0"�q�f;#.�o/c�G��_���>��H�����`���(����AF��b�$�~ny.���ebB|��]�$�j����R�˽�ycT��1���Ev�3�����4�^e0��?�59Q���OL��T+%<os�ai���{���|��n�����,1w��F�t�[$���i�~�FHL�K����x(c]N6��-[T��i�۶�?�<� &߹P���1�P�Y\�K�/��@Ʒy+�7��gxd� �bA_|��p7��%(a���VXGS:�����jy1D���<�/��R�?R�e�~̈βn���IFKB�������0�wf�H�T�����y�O�Lq�q���WW
����j$\����Kr��%�=�l�J��� 	����a�r��O�������`JM4�����1[�)⎲RA����EE��Pp&MQ7
x��:�k�\W��`�9�{�N߹���G�t/�٥���Zߕ+3��_�>z.���&�%�n�T�< �@�_��i�%.�V
�=�ՇqqU7�|pǓU\	���s���[�xr�縿���xy8��u \�v�K��1� CE�=�ؓ~��L��*��[�'d���z���5��K��.춠]+
�(V3 ����|���<T����"i�\��T��D�C�Z��|�}'�� 
��6I[a݂s�,����s��׀�7�n�����9�^15b��k5C���0�qc~���N��6�\b+z���bFw��Һ��GLA�IG�(q�����׶�q�Ў�A��A'�f��4mw(�ýF��T|�����9f\S�����/K~�Q�}G��D|{h�7�ז����5�������W?�%�|7��)N�	��_լ92pD�i�0�wT<����R�Ŗhη_�]�\�Q_��9���z�),p�͍�5n��#�!s""E�;�u�oD�e:�	{�6���V����ģ��7�9j]��Wa� �H����N�Չ����@SqG�cB}��;��Kc��uOOƇPU�r;���.jY�TO�i�L��}B �����!�!�G�NS��$�B1��K��d�Y���/�#juiVEч#�{�bG-� �r�._&L{;}�䞙�z(�)�b�t�=m_{�S4��0x�b�F�T�ʷ~��ИB�m�r�ǓbE��
���:�f8���A�Ô;nzP�<�6giX�;O�>���P����Eq�Ϳ�����{��rN�;�"e�]s��E�05�i&*��)�����\L�Fv�T߭��k$�Ё⃠�����U>XԤ�4x�a}r�}�(�$���X�T`��d�����o�!�6�R�'y��ݧht<Hx�9�����o�#^��Ժ�K�N�ȇ�_���6���ר4?�	���7�2d�'�Z�^Kg���~k����M�d��@�!R������ʈ#��)_��/�2�Gҩ%��?h,w�)U�|�ү��.���b�O��ʾ�jAM��j�"*D��7V�����)�9�)�FIM����14�%Qr��l��~G7����_%م	��X�A�����O��Џa�Um��H=v��18њ�����4NwzI���XY�WIxy�V��"��������G����mS��"n�E�I���c%����A����tc ��Q##X���H���	K�[C8!O{y"�J`W����;��~V	q�W���
��`��\�t}��f�=+���]nӉ���;wƙ	L�un����aɚw�{{� �j�X��u�A��*�1�dP���}��-�<K��p�R��1L�������Y���=���$�ü2!&z)�ѡ��
�R)v�t�q��~�'�	*-��;��Τ�G��u�(�5�ت���G�}i�	\����Z�;�K��#�	_���9�>�����'y��!��K��G���>�Q~|8�#2���� �a�`pC ����I�ݺ\�O@��0i�{�K÷��n=�H*�l���K~�CY�û2l?9����^��F���4��L�`Q˸�ғq]*�h�Gu�$��/g�j[�f�}`o��C��,Ǥ�d�5����&����)w�r��'��8���3y0"�1��W@���A��/�r0���pN���3^ω8V9^� #P|�'��sUb��dKK�=0����;k~
���f�9;����P�A�<>{p��E�c|(�I��u�!�bnQ
rW�'��@P��:&E�]�_I��$��`�a�"t*-u�u�1�b}��UB�7�;d��w֍����Gx��x`Q9dx?��RGt��[SO+�X���zGF��z@��Kr��6]C_�z�L
���R�V�+>7���
(u�c0�^ 1�;ۖ�`Y+0�3���6�d+a��� A��.���	M'7zO��Z����W ��|X<Kܬ����dt�GH^�W|�:,��j�/��v�2
I窧��m3\��jb�����S�3�%Z=n�Q�'g�tR����>�1X��45��O��pˁc8c�W{{�RXAF��_��?��v�/��7	��{%4��N��n�!i��6�X���f�����b���X���}�����7W&�,���E���t{@)�|)�f��k�o|�=��*�G�A)a��)�F�a���0��P�Y�:��e|��gwu�ro�7��Z�� n�Ŧ<�6�q��z�L~����Y?��O��m��7+x����\=
��!����庽�5��^��=�f�~�No���A����T�[��؎�5PL�ֺZ�l<cިy?������n�)���v#�]/UG0I�?h�ι8'�tkyص�\��o��v%t�����^8/p�l�Km���lT$Z�6�E}��N��`����c��A)���e@5	�59��^��V��͹qw]��V����E���P]"Rb���kX�9کGth�é�,��+���C�*7�d	��]h�v|w�ڔ�:d{��R�k��a�Qjח���LxV��L�7�ա�_U猠�#qStɥ]{���M�pf�-�,�����j#c_V�s)u��B��;���hōD����+?0���lh�F��IzND�ָj��Eb��cJ_�^����Ih�)#�1F �k]��}[zc�7�}����є�j���9(q���"߿οT��!`ˁSBN?�t�/���љG��9�
�d��]��u��Q�~�_5�U�B���p���R<� �;��
��}���'��K������~Sa�Չ�<��B捅�\��Ǘi�|�&�	�V� �@.����aΗ�-�AAK��@��E�_1��fh81K�[y&R�{bt�rS��+n�٬kTA���c�5c���-�brm#�z�n��5k7�Ԝ;|a�����#	t�&�EP�$���]Ɋ��ܢ��9qH�3<��/�bnkm�5�F�=�t�n��2����n{���{��2�:Z�*'j��B�I�>#l��?G�_�m��s��_�O�ْ��e���gew,�$����,���*�z������k�[��F�[Q����;q64g#���v�K�֤w���A\<���饅J����XN�1�IQ4EA�^����h������𞯪��J�0�u��Y^�$kI,��� P㍊B>�0Ե��:��~R=	��9w�w�h��r*�Vi�`y��%}<�!�Oܧa}c��� ���.➫�89��H&�%D7���(��� �����W���������J�4��T?���WP����Ɯ�#�I.?[u�}w�1m �?u��+F*w���ρC\f$�R������2�������2@��X��{�~Wq��s?M��D��-�2��ܾ]�U�-�oI����qD#��:2��eO����_=ff�� _k�����M�8T�d/�v�����9�_��7�V=í�&&)�Q�5{�~մw�����< S����� ���1��)���6��pd�K �#�����7��m�Q��mD�3O髋`�Q��H.�n�e����jD	S�C �{/͉�T�F*��B2�3d��rwGd����bރ�ut�tܘ����e3�6��܇���W��7�����Yੀ�&��e;��:�e�-<_�HLp��$0���3T�^�clJD&���:8e}Q�wЍ�wfǛ������r����ļ萓�_Yڪ�)� s/���mL}��m���?��$1�/+����TR���9r��^�Pr#��Sଢ଼4��g�rEȭ�"�}��p���W@�ī>aJ�P���(�XK��r�c�O��
�ع�g�����~�%�p���b�B��� ��C���u��a��Fy��M��p��7���J�p�eK�?�Ha��]����)[JR�l�W�kM�Ul?S
��,<�y�Y�w�)2���SB^�bv�'�o��&P5ܣ�6� c�~���@:���Y�0b� "5ʬr���-����9,(|WNd�<�
�%%�