��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V�h?�xrMIp*/�p�xV��h��K����.��V�����@�u��b7VK	�>iR)�~�
}�l�	��I�T9�D� �1]qU��JP�� #.E)v2z���zS�P�w	�O)NŐ�o�7���g��_���f0�L�l;E�n�z����g��\[�,\h5+]8>)܎9��
��#ɝ���gK��ͪݝ�J[�o{5Ui�g���^�H\�����<��h���Y7z�{|�0����d6Xo H��Aڈ�����!����f��"L�1s����{�/S�O��.�m���5�yAaC�g4w��x�tu�4�ݿO1��tb`�uʐ�,�l��J�~;Iuz�m ��A��� �;�9ĖC����c��*�P3
@,Pj��������;M���R9�?���r���m΄'m�}��������@�gf�ڤ�5�؃A�6K�YmsH
����*��.&�"�"���b�b	�1��gB~����7I3�JY� �]�.������@�b^?yۣ�NeJ7o,������#/���J����q���vxK>�j����0� �o�ߪ
`�7h[
�y��,�MD@'�^����#>�Zt�q��Xf�3�yME��jI�2:�0Ƨ��=s$#Q��=�瓂Ol���?.&D7c�3r�e�[�s� qbQc5�S��F���4�Wn���E
B@x-$�J��Kx�ŚoqZ�{2X�r�	�p�RO�#���n}�ڧ�-%h�?Y�3�C	����ˈn����B�d�PDX��]�
������s��a!��p�Ǯ�
�� 4�����c�d�Vߑ�����
�6�E��ݛ&����`�`����>W��z�-��c!b�RLٯ�s���R�ǚ⦎U{��C���V�%�<ش�?�3�n�&�B~��$2ػU�
h��`E�ƨ��!�$��aG��Dv����OU�S�]�.��Ŋ���Ą�*O�3&/H��YʓR�K}.�����VM�c����u��$<$X5W�su��܆���{:���#>غ�!2����}������'Vvᇏ�=oeZ�l�ۦ�Z�{�.�"��� Z����'\a��h���`��#q�N��r������%�b.���aɩ��~���Q��;U��߱�9��Zj�5\���������@�F��t��"�QzWl�f�� �7y���'r�A6!@٫KxE���r^�l/@m�x�r��-���o�����R�����H�ۅc�\�B���tM-��>�m���̜x u�3��
�w9�VԦ9���m˶<I�OHc�o>Id�w3j��rڴ
cw�d����K�з���#�@��t��
�HI��hܙ��Dm��XV�L�,#��j�7�Kt��>�	%� q�����&���x��}>kRb�G���(���I���SW(Kݳ��QRɓ��9�<t1��(F��#���e�����@|6���Z�G���:���ՎՅ.^�̬ܩ�����ն ȡ�
����8PsD*�\5󞖕�[k*�{�ƀ�u��86�w��	�W���(,�n�k�E���N�>
\ec��;�������+�m`M%��x�k�����9��Bd3��z��Nݍ�ju9DO+-�0t�=Ke9���ѓ��H�)c�솞+0DZ��8c���ɟ����
�ҵ��wL%���fpɶKsjJ���&�ۅ,�/;���ք��J�F���,��"{`SeN>Ƶ#k����.Qկ������ָdIȅ�N8E-3ԝ�B��ݻ�T��x3�i��!��x��< ��]w����L�occN�	&�$b���*̭�$ԏ�c�cO�7���b��ӣ�W�@�5�Ӡi�rǘi�Es��)���S��wi�	��bN�p�G'�Ͼ��drt;̀�e�n$���(��^����#̿�b4�}���}���L��<��Z�i�֙1̃S8��J�Z��"�r�B��&����
��4a����w$;'�����e���N��p'�]Ɩ�6���-L�� ��C��t���ƨ�9¾�%i�a�fH�X��.%��A��XU1	��KK��y�(��_כ�h�[)-[�����4�J��U�ο��/�?.s�B>bF;X8X{c�2�pW��
����S�w��Ǯ��o�&�+�Д�.מ���1JdP�o�a���佮�1��Al(=���F��ei
K�f�&��~��c�5$6X���R�V�q��-��8)ƿ�m�}��.��v~x��#Wh���˚`6uz��D�� �a��)�!)IP�+��Ҙe�����N�8XH��MJ�r^Z�����рűq�no�
{�*7iNKdAgt~R�/6�Z�+-p���эojK��V��y^�s0ԕ���A�b�1�f:\�퇣�6�0A�AD��e�"$UF+������_(�	���h�<��l\Z
�����
�: W�)�"�r�E�K7�n/*q���z>A��u�fdL�����zI��9ៅI�aZ������y��eMM>�s
�{9BEGW�����z̾�l����*�e톰�wD�n������0@�t0g�J��ӗ���.�ḑ�d�Dg&N?�g�^�`8�{EʠL�#��6�`��d]���Nx�jw��P@0���Xe���7Ym���63��?�[�`֞k��!��]�Qo��NCk��患E��";�ٻ�y|k�;J��� ���ʣ�+��[�{�����Q��^��}�&oޱ�?�q�ف���>�T��4b7�E�Y?��7h$�9�	�zK��`CL4a���T��"8��?��%O_>��:���}���ǿ��*�ً�`�NȬ��z���4�S�ն;�C�F"jJ���IƔQk�.}�Ap!�*��U�P�!�yc 0����;|7NC\r�����5�zn�P�/H=��#ABs�YB7��o�_�wRv�m�6���H���7{ed=3,5o����[�:��|�?�\����L|�#�^%�M��Tk)�����h*��i��s�b9�a
���*����J��yr�dU&&�����F.L[��~�k-�����ѐ�ě����\��,�Ħ�H8�O9WJ��x�<�l)�E�#5�~��h�i�n����@E�V�b�`j�'���Е�	�o���&��R�`V}w7�|����̊���Aa�:e���jN��T1ϫ���k�$�=M �o���I���� 6JIg7�6�3�>H��
7�͖Y�)�vѝ� �l�n�j�u���W��_'8RZ��A�g�V���g�WX?�qe[�S*S��O�����&�c��+������w_�_Bm�"�*�
���Z���J�G¼��?�l�)�����j����ߕ�����K����$[�R3NA�I�xbSNIU7��^?�S��AX6�x�j��5l�HҼ��/H��C�g��� 9Y!�}h��&$�N��8�V-�ͶG�-��pdcV��Ut0��L�X��*3�%6?ⲥ\~��	�p�X��'�����^<o�P�q����]I��b_A�k�}�"_��򇡡�ᗅF	�Yf$o=�� ϗ��V^d��I`�Z�Q�i��'��B���a�����9�;�����>����GX��^cV�pc�ݯ�H'A]:^�RJ#��0s�� ��`��o��]��"���$�@d�˱����XRB�+ �?�д�R�%�9�HS�˛欭��=��*H�C3�"�7�r`S��
[��<6�P�s�����t�OAM�i�gdƔIT=�3/桄jZ{�P�_��%�mĂ���0s���l�{�
�yE�,�IϨ\��W�\W�n(��n�Ƥ��y��I�fծ�-���ƙ�v��j�8���CM�B7��t��.�&
��+,(\��q�@��- �A��?�)��J�m�F�Y�CsP���!�&%@/����}0-~P	�	5u��%�v���J�s��ٍ�*�K||�fkH�WAI�p��bZ��qT"�����hO�r'�A�e
S_Sӗ�( �Q�>�a[�!��[��P����yE���s_9����1�5���z,�fΗ�����;�D�L/p�u˼���&��ζ���3x�Y���/k�'=��%�>�7��u(q��5 �O��<2���#�5����7����ܥߺ�;��m�z����X ��1{�ŵ!��"F�1�k�	2�ݹ���k0�n��N�BP��#��C'{����l�2h=/豿3�""�Ĳ�[qD����െ��#���]��,ahz�{���e�=�׉�D �7` 4� e���ET0���P�aV�\A~�KqGz1��hs?`N :g����1��a@��$��u�#�d���hnV�w.ܹRx���z@?��t��v�λr+|�*n=Vw�����+G��;,��:'nG�l>چG��~��n�E�3�O���{W��z�IG�1�mz��8������g��rK�S�7,���v�l��
��@n�_����Kg�ɛO
��G{��Z)p��e��;��D�Cc��l�E/`����$��������ҡc%������iv���O�2����F�X)��۾���v��v;&�=}(�?��� ̣o^q��8+`���*�Z�4:��+���_)J���rf}��Ċ��5�RjX�V����͈�z�z�$�J�Tu:�N��$(g4ٔ���N��|������(����r&��2J��$$�>F�\OB.4@��M$�[yS�8l쏎��d���D�y���VjI���w���u= M°q��H�������K�"�,���ڭb�}j(�����v�X����%��^xd6 8����$��@��l�j���)%�$���V�%�p}M�P�S��'��ux	�5�i��`�f�"�-�(1�A ,
��
�+kEB�NݩB�;s"P��_&�4�B䗏�����z��^N��'�HhPsl�L�-ݝ����F���S����ZZs2F
%�/U����9��D\'�4�� ���faNo?O�TS\�A4 r��+-��o�� ��=� �	��|E�I6��C�髸9�'&E�7Rg)3��q4n�g)����hN�3�Ebv�1�S��c��F�8�f�J�"�ŝ��c��!�����Սz8pLkQ�6�h�6�+�D 4�ӟ(s��4���:��o���WbZ[�H�� /��8;%i&���*�~瞉��L��E��I�������ֵs�����y��ʦMv��3�KR��C�]6�&q�dʡh���褁9���R��@��u�,*�
NƟ�T�_VzR��֦�W+��=@��ZF���!$�Lm�6�[oa`B�|ޑ���[U�G�{��*h���m��.���2/�����B�����Do�����Q<?���A���35��"�zlŽ����U3PM�8��->�p��.2|�j�L��%�iW��(*䲆�����P~:#�J`T�7W��m�
Dԩ����E+0����:����3�����Kj�j��n.�̂S���z��pjP����E(f9���TR��#?��b�5w��K�\��X�S�[�9�{�Y$O�Sbg �%����$�a��W9}*�(nk�s�jJ#�u[&!O�q4hS=�.���sy�Ƨ�޹�kjdDs"]h�ǖ��^�lK��u+슰�S�Y����r�8����3�m%
�4�*X��xz��"��m(�T�R�l�Z0@�ӟ��L�|�R<-�Q�#UXq2�KjƯ�*�O��-��3)��A����o����u�#�Z�洠Y��~�f��������v�~��Fp*�
	Q�96K�?���E|o0=�DٕP��^�H�)��zWx�M�k�kb"��Z���B4ב7�O�{��,�ѷC��"	�v���K�x�|�k���i��^��r�c�J�;9�88��1������$	u6S-cb�2I�V|5R��/�Qb�*Ui�&݄���`~���S6���EoՉ������<=���4�:����͌5ƀ���K��u��.F@���47�c�O��f�i#��d[n{��}���x,����[�&3qH{$�ӏ��W�����t����ԧ��S�XH�#̗���;�D�� �#ȍ�Ku~�C!��N���hv)i�%�XJ� ��(�+���/��7�2���{�/�或������~�{ݡ(����%�{��"��y���v'���si�>&����أ|g��7K�C�4��z��[ON�{�U�����NR��^�	�s!aЈ,��"���5�ۓUDOdP��`FH�0�o��T�׀�v/{���E�c�*�!�\&N���N���m��7�\;MG �m�j�QǴ�D����|���@�(���@-�T捭�Z���9w����*�lLȁ5�S�S�Cz�,�G�9-FO�Mouؠj
���v�A�>*��؟.쎱�,���^m!�קhG��E��6������*��yc�*��p ?T�A2�Z3��2���"�5�wK�lEx��˨Eؔ+L�'������FN5E2�7I��_
��rq�_�;{�:���E���/D���y� �l鞲��H0�c���4jp	!S�a~��e9Ơ��y��$5n�,tR>t�$#k������l�Fȫⵅ�b��s��q�V������{��a�5T�	h���h�MF��9k%������t�u�A?��Û�~�(���p��1�"����[�:����HH&�*�������T�"�7���}�L�Pd�5�U�3ږ�	��E	UD�|Iw�ĐPK܋��T屆�֒�>,ee)_��}~뭂��^�\{$�&~G8��6����������8sL�"�0�[p>��ʟP?��)݄v�i�h!T�x2������ªC����0�����X6� ud���&�w1�m3�21��Q��}<���5�i�Gd�V7�@Z�) �$Ze(eڂaoêh��l�"������Q~��f�+ӕ��<��&Þk����Pi�����:�1�q��H��WG<��Y�d1�gK'zMC�gK��HՇ�����]��^����g\Y�2[���T��u��rq ��̠����5vslU6���i�߿��]�ў,�_.��	�}������MZ�eRn�_�@=텫R� �M��i�O�(�A���ܖ������pM[V%Txtw�ׄ�M�A��VL���u�J��$R-ĉG�a��}̷9BX���{2�D%�ݡf�L����D����5A��q���H�¹,�O�m�k��}^	}���BN�����W���l�1���=1G���F�VaX=�mEQ��X(C�($M�-���"��ʤ ���Vc�(�3
<�����7K5��$K;ݔ����?���9	#�7��9�o @���xu�P���6_��)��lD��S`�!�H	��(~.$�K�k��@]n�{�=�{�а�!%c��>�^�>(=@�U{�>��˫��b��U�\�>���P)(��hj�9ÑV���z�⋍��V�*f
d`��J����sr�"7�7~rt�`=�����|
Q]�	�Y׋�t�z>=5��ԥ%sg�oi�ֲ)�����n�Yg��R9�DGiY�Yj��_�Q�!�+~@� ��ϩ<R�'uG(W�aY�Ҧ�(-X��)ĸU�w{9CZw���R�����a��}&���,~�U�p�x�	祣R�I<�=�N����K{��iI �Ϯ&���v)L�'�8�/N���ty������*�5�V��`�I;��T���#�S��ë��-��~P��I�c�T9���5����~e��H:�=�iږ��ض�%8�U����p �8���5^M��Y��</,'�Hܶ�Ǹ��$�����*��!���(<g`�N������p�ڛ̯{j����Ƞ	�����`oo�B�^J�E��M��U;������\���u�(u�3�\�̕��A�i.�	 �;.��<�r��z����?h�{��:@H��d�/`��8;闟���Us}{��	׊�������-'��J� �L��
|-��	x�E�!��cd�sG�'l�gzR��&>�����D2�O&��=Z.�Z��� q�+u��8�u�W����������訇}#Ɔ�D\+@X�>�~�N\� ��mIB+�0x���z�_�^����ď��ʀ�'Mf����Ǹ
�b�4F�5�}�B����d$�h����,^��Y�������k������,#ώ����Mi�v��ȡŠu����n�rA��Z�%�&���%�%�b_!gܲH]�1l�<��a���ҏ����<���Q�{3�3Ȣ%5;�F[��#]v3K\$�o-�U�&Bli��F����'8���I��C����l����C��^��$Ew�W��'{�`a�U�74������Y�7z�"�;i��ȋ����BlT��CН�6R:l���?�X2!���yA�3�㩱&d,'"�Sf��̳R�����OQ��d%��c}��`�@�ϊ/��|��-�\�Z���)}��u�`��%�ɐ����$��+a�E�E,���������h�f�61O���n�8lC닱VX^C|����X��=����!�����c�ݪζR�>Ю��!U�ڌ�
c������OQ$MA�8D��W!G-݆�H~e1S0C���A��#@b�{�����{VE!^�Oed1����Xp���)�L�\�I�fp�z[�U)�f�I�GC|��h'�P�)k�0��W������w���T}������-L�(�MI���2BR&��߷��H��^
깩O��Ō�ǻ�r�=�^�Uc��3ѨV�4ѭ�ӌ�Ա��Zt�q�XfP�¹�z�_���v���6XA�U�r��Ei�%��jT�'�8��1��-�;y�˛����뎟�Y�8�̒ �3�%-�M-Y�����%hv;��i����`8#Y�HY�27���n��h��#��"�����6��� w��xb|���6nnyq8G n�I�x$^�ws��D9)��`1L�1�6�E\@@J�'a�օ�)�(Gx�dM���|�!��C�b��(2�hF@A�ݺFe�R����C��nU$���t���G���cn�s{��@��5
.j`����MH,n��"�BHu��g��]�/��0� i>D�r���{n�mZ�bm�a����d���ƶD<�=	1�g��)���{l�i�b�{iT��*Ä@/$�t��Tse��E=Yz���z��%�`�U�5Ve�go�_~�tm�!c���8��F�RQ����m��C�$�)����5X��
�����9�\��P �,ج���j�d��Uq&���'�x	��y����|��ؑf*Z�\��'a
��f/�$�4݇M�tOǧz.�
��&^F4X(��s�^8?sZD����M��>��ۗy��zR!�Rn|��>��V�7�Q��};s\��[�HgZ3���w��F��w�o+&�ť<�������K�T`��H�]�YG
���lS�=�Z>�9����V���J�f�� /��_�����a�5��)Ј��A�JP�������:�pȼ�A����~A7���~W�J�O'�:3�V�~V6�>��8�7a�L�֓��6P`b;k��;&*��C�4-�ei��~T��64��8{��v7�j�5�'�m�2\�Lנ���.�(g,��vy4 'F2��e�4	��`��2�y��D[9pk�S�)��@����0q�et��=��I�;�D"Hw!cRR�<��bڌ�$�W#�������H��|�9�v�>���Tqi�;�Pr)\��PjA����tz$�)7q�AS�Nϼ�M�x�:j/s��g8)כм�LRZ�6���ë�a���+�oS\�z�H��ɚ��ƞ���v�{ ȹ�:���|+�3]�E�=���&��k̺��8m��^�UNˣ�NyuW���* ���hr:��\9-��2*��7�%T�zn���t�A1
È$�����萵.�:BM�n����/�&�%w����A�t>ŉ���bN�Ās����}���6��v���w������:8��zx�f���-{�6MQ�H�+���*˒MA�TBva�P���\=6�"�k�%:��/��[����5o�N��AFq�+"q����Y�("I��`���攩?8`�[m^����������6S���W��z��g�M(tST��Y������@���{�'"(Q��Bars�w ����u���q;�tSUY�cFL�#lZe�N�I�]*��
#��������P�c�x��%97��w_5�/�y�6#�)T���\�¤�D���5���M'�`��F�T4�ntZ"�v	�p�Q�c}�PN��$:�j
��sU�|$p�v��nV��q�8V��w�#�w�:��(�	/7¥��9ǃ��-��Bƒ��{"-	�NJr�#a����2�gU��Z�����;a�+�$I2�Y�&3�����;�����16���+��H�T�̟�����������o$	��弾����ݼA��J/��P|d�/����k"�N�>�}ż�%p��[M�)Ga�&�����ր#�)�ִ����BtQ����>���Yq��<�~sx�?|�)b�� ����D+ա���R7(n���US����������Ŋ/�M�[>�^�n�o�qʅ�Bzq�K��h�������暏�UЦ��d��sџ_>"��bF#73�w�����1A/�D#���r%4�a	��7��:@]  <q� �^.57�9�X�߭�����zZ
G;o�X�J����+���[,d��SA6b;����h��|�!/��T'D6�U{m��==0�8bF��4A�<���5�1�}�V5e䜞 ����^?�'+��Ac�s���/�?q��1Wt;��*�T-��r�6è�|~���QX.����`g٢��h������p��N�S�5���e�8`"N?{Ǎ�ʟ��&�Z�J_1_7a�*��n�a9ϛ��ʒ}?��_�jec� "u+-�9�������g�VFO�q����R�I#�����<���Tٱk�`e��
��7N��'.fA�z�3��3��F^IP�&ʻ���P���D>�Կx�WZ$Jɔ���d�N*쮇�܊KE�z��|nv�+���DUiü�Z��� ��[�%�;���*z�+:�{���$JnǪ��NH ��h�E��OA.����.�{�n �� �BC��LJw�Z� Ė�����#r��*��%�D4*�5c��#u3O��Δ�7:�<��y��_M�4��aA_���;VҀʌ6�+��|�#t�!#bX��wZKD��4�?���B��`�����N·�x������nS�F��~yH&�ˊE��W����	�c�ɺ�>b��%nߣ� }_^�K`�A�$h��������u����r]���l
H�_���Tv�5cX��fkHG7�H%���H��]r!^�P��^��x*�ac�j�S`��}I�o���*����Z�Ƙ�9;'GTc��"$"R<�a}u��x���Z�:E6uk@IA���k�
($c�L�;���Z������߇�A9 ��#��D�*�Qqt7������{ةɹ����,�b���1��r.�#��N=En�|�����!v&�ߨy����m6�6~kJ�?M�B�[w�������\-ӿ{䔱�w�WP��3�� ���� 7��}����ML��})F9gVRP.Y��g����
_�J|�2��檁CȓĬ�O<2q���b���U�v�z@��'���f�a�5Ni�<��?���?錃R�O�b�v��M��k������y�.��mPGB���*�f4��i���Btῴ����6�W*�(r��$?y;��,l	1�s�N7��cn�J7��61(�0��6��
����.)
+�#�Pp����1�t�G9�x#7mɖ�Θhg��X�j�OY~:ǆ���&���&cճVS�k,�?���j�w��C���E�݁�1��%��ã�$�n��:`-]��	�0�RaB�|��{ջg{��ޏ0��9�O�I3�p��Rz����}��˽�E'�K]���^x�]�hMW�1���Bk�M�����F�6��}]��hx�r���[C.�PQ�	
#�q���=},i�+��itl� x]qd�
��z/ä� ��x)do�K,wX΂D����}y�dV��R�`F<��s���m譧�hsY�?VQ˪d�G�T��Q�@��ͯ ��@<0�.x?�j���לP�1jl�dC|�ƕ�t��	�:����.��Q�7��?	�z��:���{�[D#ƀ=P|�����#�������-���:楛���>��*QĽHA�!�h������-��
+h\��Rs��p�3��X.��b��#�ZJ߫����s��UЬp�܁�:̮8�Fc@�ջ���nn,RIfj������ �c��Xn�O��f�,ݽ�#��/�I���#g���_�m ������	;��6hl���1ƒ�I"��C����$]��η��z'V�iC�W� ��	dU�������8T3��ەH���)�2[û��A�n���f?z51"VDs���3؞��+����Z�&���ǜh7=��� i���Mh�~>e����8g�F��q��8k�l���-uF<?aB��dd1�i9c��o!x����$�&��\�� ��Әg��]d�msh�R��\n���`�	
�&{SwNg&m}��L�B�)��<i��F�ڢ��-~=�~��W�e��d�J�D���DU��|s�W
��*%X���<H4���w(��`��	��[8�;����#�2#��Ѭu����n�:�����N�֍Lˌoь'�J㭖!��i#i��jd��/���xa$qQ�v�)�;=��<A{L�j�CA���ve��S��o7��/�`Þ1%p���Z��K@�fa�]��r6�@����;]�` Tli���(�Z������bFd�N�M�����f!���,q������_]�U_?"b�'bR�����-�ϸ�İg\�V�$ѵ#�i$�EOZ�D� �^�z�=?.��*�\�$��>_g�d!��T�]��l��[?��+�҇���=�V~9.9��)N�P��+�ZIL}�{��sk�i�ŌNg[��)���yR��&��!Ua��:�� _�7���`l��̕�q�`�L�f�I|��pe�e P��,-frW]��\�\�t�;��J��ef�A����&bmM�LzQ24�xB7 ^�;�Ⱥw���}9A6�H�@Y��m��U0�K���M1͕��3!_�S;NƝ��j|MRA��~�|>���i[?dkZŧ����%�B����D9/d
�P^Z�Z�Ѩ�[��J���/���<[�W%�*�Ig�C9}v3xzB�+}��.���~>��1�D9V��l)��8�qq�W����o�P���"��g�3��?��b����W�	�wHP�����������9m�y�@��j�9�X*3���LC	A(-(���!�����b[�ʫ[�d���8b�8�Hto�:�C0d>ܱ}��O)��+��Ab�K��ulg���fÒ�0&��K�O�u2�B}��S�exf�#s��E�� 	��	�g@�I�`d�k�V��ۃ6����<}�� 40h��G�Z, ,s�2�ո�NG�&�(Wo����Ä�*���d�A�o\��V�֑�⫪����S�0��������Qƨ����$fJt��P(������p�����ܲ$dw��� �c`|��u�Mм��v0���n�p+`l�lc�%������� F���cB��VB�����)�4Q������=����	���(1��q��#�K�u��r�S}Qj6x�ہ�.�G���Dg�8�\�R���f��͸;��ɴm�PՈ��Vn/zwjE{�eΎj�UD���
*�d�$����x��ފ�O�����$��|۾�͆�0���@N��ڿ �1'�H`�8<x�p���|f���Q�oW9��!oI�aY7�>�ׅR��Q$�'J
�<-��� ޔGk�z6]�wk�'9��-����f��4<����h1qtX����V2s�t_%T�0�� ^��V�U'G�)|��x��.
�ar���Ժ��e�Yw<	�*)6�@����=Tq���0��u���OT���v�L��>y[l�ܢ�>gK\���eD�=�ÌR�,(��L�e�b��uC�BLD�C�@ţk�AI&}�hT6aR� �!��:����g�>d�簯�m�u�a����~26� �����쨮B��7C���e��C �&}�� �E�a�u�@�x#�5���˵�qG�\8��E9Qw�݄bb.�QT�d��S�,�V��ژ:���+H`x<���J!��=�Қ� �ta����z�t�ЪIGZi�����84��NO�`z�*���t�G�MW�&<��΃��O:c����Ɂ�*V�SX�u�E�.��<�lng�r�a��ic��'�e���+�e������Ԧ���Ҷ�x���B{�8`�"�F��Uo�(�>���֭􄅁�1�h��`y���|�ԓ�+�Wf�'���t] ���L�%�yw����襦o'�A���N\����"�>��)~Ƅ������cL&�Ϲ�
>���<�l�g���^Ꭴ���L+'�wԺ^�ǘg����j�?�����s�~^0���&�[���uk����8}��ln^.A����qW�W.�Q7/H#��0��c�&m=P��͢1�Iaڶ�e����`ɨl��l����Wɲ�{q�O>��n���&�@��/�<V�����y�9d�!S�y��6r���
�*�Bh+�y�z$�+s!�j�?8�n�L�D�q<ܖ����X�ht���ΗU��` 6��A9t�$e:�q�U�y�.�Wo8�ߵ��}�I�S'\J�L��'�
�)`�·�p+
���F/���(i��t���������ex