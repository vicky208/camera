��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:��r	��a������8:`��*ߋ$	��L�<Wr״`��Fao����kt
4A�tX�X�􊎠y�Z�Vȗ�di�|�_hpP�<~3��G��~
��t�0��}�]wm��=�i��皜f�+��!���ۓ�>1~%N*��߂,ͪ���*��hN��u��.����V��U�e��ws
�W�!P�' D����*��<��d�R�i��]I�򗏴\_gl
�d�#���Ivv�Ì��
���w�z!5�,��L��주	�rF��!�]G�p�`���J����>A�b5=_j�pA3ƒp}�V�$�!�1]Զ�Re��kĜp_� �c�C~��"�+s��9��p&`������ן�y^�i;Pc��	�ns!> :��[����Q�|[��Ʒ��:��A�cnqQ�Zl�.�F[�qr�Sj���yܨ��X��.׎��u>z��ˉ�ʼc+�/��P�q^;�2�^����4aE6�n0sWЗK���X���)��3GI�[wk\r����č8��	&�N�#����~&�����g�XR%�����2�kO�'�������~b�n�E�wq����g>����`Ft��htl��}]�����-ML`0Ϩ6������m�w+�+��N�t<��v�专w�{�T�EY�'��۶�Ī�y�U9��X�������L�C)�`#Gl�9$�OX�J���'_�0�$�,����jw�VK"G�Ne����,��v�����NqV�Α�^}<�/^$��
?�b0����7M?�'�Ա� ��*�\�OP��S���_z*+�X���W�����kfn-��^���iT�:Ma���BH4glJlz�Ҋ)���(C����9�պ����q�����r��� �8���xV,�q��[j���͉��0�>��p��&����0x����L/��DO�X���������z��J%W�"�I耐��t2�Lp�e��zL���D+��%|'��Y��	D��C=�-+���vR�e�d.I
��K��$�s �Q�����*Ʋ�����Mh��Έ�y'�S���Z�|#��8�V�{���"X�4�ܸ�����tÐ�Z���b�Ai�������#�e� +����p�h���?��EC,u�Q�xI?*��;���*��-j��e�(�7O8 ��9��21�WqY�^�{��P� ߐ�����a��L)�@WUk���"�A�[�"�[�XA�D�\�L�ڻ啫�ބ���o]�Y��JI-�Ǿ�-*����-w�w����ɱM��a����`�"��;dz��z�M这�^m2*[��n��X�#��?dJ�S/���ֻ�x�ѡR������f���߿�@N�#?�ѱA��(2h��'÷���3C�ŭ.���D����Uҝ��#�_b�����Q��>�L\��)�׃u��2P'7G�k���&��ǀ^-)d�m�w��7�J���܅bC�uҥ�0"�NE������B*M{$����Zl2Ց=[��4��a#���5����A��mm�E��rLE��VdYn=\�E)Z�?��o��#��S����^-H���1��|e���s���Z�MMr�	e�P����Cy`�Gl� ?i|�����lv�\�\��Y�w7OBnJ��/#x���g7P�8�l�c-��_���H�)���	���=��8	���(מ2�<�]V�3����哱�0��y2�^A�����g��}�WΕq/Q2pv���B��ߍ(��t&`�!�\^ꖭ٫��"�Z0T[ ������[���!0�
&���g�Sh��V���Xz�x����xp�K�/L�Wٳ���&�^O/65`g����C���HY���A�J2ԩ����h+�	Z��ǣ0�X��˪�\�K~�4�ȂS@�E=Vs����o�^]���x�ߟ[w���UP���0/��C/�M%5��Ђ�u};�$��w?�e�Ht�Q�]�L[X����~�h@�oq�ݮ�1��({O#�LvJ/ ?��-����<��Dc����t�%ִm���[�t�����xC�JDs�9�͒���p�\��X���\�h���D�j���;[9n��Q�������P�x�n�~?�U�}~���p-��^�� U2�*ｼ�@"a�޽��G����r�����ߦ�iWn�W����&�v�\D,��� c��v+h����}�V��M�{�e5����F7�Oz����=�����@�I˻cfk��xѬ�s�Z�Z�*y�$ZtwK�2��'|�zr�҇��		ZG52	��z��Tf�P��{[+���*S��n���	9,�VU���[����m�z��p,]����x,q7訑�M�'A(���e���hȫo�Ytc�_Q���\�y̥�:l'%L
b^s6�ܧ��������/�t�.���d9�Qn�X��+~�����\�.�)&]@�i��i(�a$ҏ���fnm�u�Бv�Y�{��IAa��m/�<ul�v� ��_JH�=~���éb��t��X1� ޽�[�+JU�����2_y��~z��c-�RsI��d'��jL__�b˲���9�(@�QA
;�+V)>�[a�9�ⓟ�h�x�a��a�1 �b�(��g�B6t�᭽�`<�t��V�An�R'���vǓ�0��.�����"-�@9 �V�*����<���Os���RɈxR���3�3EV(�Я	�~�$2ƢF��ؓ��z���7�*]+֓$��(��vc8�����������m�l�Ք_?�2}�u����� ,��p*5�퐉cB�\ݐ���lH8d��|scb�N=���T���7�[�G++��e�u�4jc�{��KS�-E��[��h��������%1�E��"���f�YV8^�B�Ag����!.�PN�KX�F��{����r�������yYZsF"�{�߭ى��!��4�,I]\h�K8?��!7�8@:���Ϲ!�?�V���*G	�Ȅ��5��0]`N�K�������oPVUnF�`i��AIю�~�{��1^�ޖQ)��)B
�f�j�ݖ������Z`(§@����:qԟ�����_ 8����|�Of���j	���r}�����B��6f͎������>�0�ϑa˜t?o���S/M�8�d�1�
Hg�G�<��R�l�3z�8��o�A��b����X(���Fmۈf]��Y��&&�.�;�=w���k}��t
�ߠvx��e�wJ��o��s����u�����_[f{n�UB�i��5xP��K�=N�-��K�/%a���q��Ͻ�����q���c1��(�IGOg�
Q���vƘQu����h����-fc��1��3N524E��+��j��/��@��ʊp��*V��@l�Nso��<�
΀0~���n����'`������`�2��Q$��L�^5-�'n{����aa[�[Xﷇf7��t���Kd8;ηvX�\8巿��^��G\���&w��ν9�ծr��|�Y/�k=��3��N)V׈�[us��o�L���c-����G��B�I�����}���)�u���h�ͥ�uZ������2β:����ϊ�ߤ����q�-�-l�[Ð�2�k���L�`�i-t�l;�VҸ�S[&��f�>7��gψ�HL
`�/#�6uV+����������Z-����
�`��`F/�I�����f|�9M���gl�I��}Xb��'���9]�;)}��8K2w�.=���Jo3�u��TIB6�}st�a��~Īl���:qȯx�ۅ
ň2B럔L�wLkD7�������ײ-V�`1���^IW�5���o��G�Qh0��2�L!U�b�C�r��]�(�O<����" -M@�H�?i�����i���+�j�m����Ic�3�R��v����5D��o�yu�8XX�o����@\��7��i�*s3vs��Dw�{^��Pp������ �v��ϰ57��m�H0����! {#O<���ԟ�����zc�;�섃o-f�$.��}I�JUQS�]�`w��	���\*t���I�/�~�R�H���*Ma�L�����<|3�>�4E�.��yHm+���o�����9j@���(��L�atBQΪGv��� 8�s��٣S6nA��oC$u�uޟE���q�(�/�M�2��4�Hc�g�i���	�@h��	.̾��1�Ð���1)@�O��~Wc��9.y���������2�)c��w��"��1��<�j�]�l�^۹�_��xdL҅֜����ؼنZ��p����+q��N)�
x�;��CY(mh�=o��/IO�����<����~����
)9[�?:�������Lh.�V�T�9��$��NȥC�F l�p�Q������$���H��TmP>�e�+οWR_2��<�W��f�l<I�¾Z�dw:�}�Ԇ�b�����H��%���[ >$���?�H��9{�!3;��P��G�I��h�\�]}*0���~��s��1)���F ��.d�h��v�sn�6\���>�{�˔���:�,l�<j�eu�z(}�� On�F��d�u$mR��Bʸ[cNyM(8Ҙ5�*��pM�:ԛ�]���cJ������}X�Գ%�T-�yv� q�ƺ�?F�nO����y���N�Hm-��M�ƄNng��1<L@�E��%�ҧs��{��*mv���2Q�P��P�G4��p�O>�]G�>�e�;^�"�:W�k��iv�e����V#�^�)�L/�!��6%Sǡ���
V=�tb��i���&�l8ßH���*d���=hg�h���;b�Z��f��s�L�e����\���f�35�$�"�$?�p
��<��t)��j�(x�/ɍ��T��|�w��u�&22��r�K�.���q���v��o}��*�ڳK�\�6M�r]c��sE�qq0������K�5���P�9�{��f:��V�9w�1~�,�B��#�\��n7;zvV�J���^��d9SV�5�������V�L��
�.1�*M�(�6��}�*Eb��,�3�d��󨊃	"׃e������;�����u �^O�R��.n;9YZ�D�%a�֐�V%�Ѕ��<�����^��r�Y��u_�r�\���}����9]�R���@DXMj����?H�n������_�Ѧ=A�1�z�|�*P=��.1�ڐ�0��������b�@֚�&8����s�Z�L)�\]���+"�V�o��W������x8�so�e���Nk�Xʖ�[2��%#f�!�9\�^Z�@���\i����ia�[�%���"��n�C�)(&2,yF����T&w���"(a��YS*&%�yȿn�D
�{9��b��HWpn^g�O

"��A
����"ȀȦ��;��E�3��NE��ѭ��Y5��?1�S$�IR�2/Wգ(�e䄟�c�g(� l�v�������\mB~��3=���t�KD��iӛJ8rC�g���x����5�����'�.z4=�*=QMWbC�nu
��xc-��{ᕢd3��k�[�_.=�j�ΊU�AQ�o�P�%�Lȏ;`�AY�:�((2�,-=��7��z�)"�������,z��@fZ���L��QV\�����0��P4�Mk��mZ�<
����O-n ���{Lv�#��Ō~�k�H:IaG���W-�)^���G}��d�JY��V��h����2�:6� 4�n��~j�|���1�G�w�$7� ���(j6t�X�q��cǼZl-!��PA��2�|b�A�H�t*`?�{Oу�ɻ�_��}S)f$mO�r�?�H��� �2��״�D-ndۇ���s	 L4J�t֧M(�Z�f{��������,x܋x�����,XRд��ú�V���0���uT!�R-h4����(TȁO ��i��~���kD�[[7���㠘*\��ɘb��(��`��D4��(w�GD&��Ϊ�u�>�Mq%z0�zci��x�k` ^���-G*r�E��3QPgIh��]��-��Vg�r ��@r'F��_�[��I��*�~wZbD�̅)s��l�Lx�ѓ�m�p�$�ù$�V�cb�N��2�T0�,
�r�Zv�ͤ^/�l(�-M;@Yg�.� mB� �Y�b�칪,UA �OWj���\p����U�m� k�}�-��UF�/���Dqi����Ĩ��=�wh�A�e�f
z�������gN�T�"(�T����ID4�0`4�^wV$}���	��1$�����B���\}������^��b�l68�#���6�";�N?��(ٮ�#ȩ�	���m#"�wNp�D�nd�����y��0��ڧkA�x�=��q���
�EQxV�VD���-� �lEI3�Y&��{!�>V-�s�kS�Y��h��_H�*�t��$�e���7��v�2�(oA�Y������S���)��psy���y���I�r���D��ǠU�]X¢�_[E�n�}�-���;���O焚��M:�r%t_I�54�p�'u�ܯ)�y���!�Ni-�������S�����S'T+�]6X1��&�(|��N+��-w  ��::�d2���"�7&�	���`Y��_Fiޥ ����7� ��\Y��a�ʿ �qj��AV��a!�EF��1)m��b�yJ>Sg���)B�g=�¥a�M2e��:�o��?��	c-��2f��X�M�;�VuL�8br���O�QU��70�p�:X(�����"o��nߢ=�\ �.'
~�~0����d�ZȎ�뽻;�3]������b�A�F3�e��pB噉�g�]���/�5:M�

}u6e��5-]u.qo� ^�-*�I�����<Ɓ�Ř�g#eʯ*Ê�.&jV��8M�u�2&�`Mr��Й�03��!��<�\�5E��zp�Tw���Ff>�Sr~lxܖsXװ����J⫌?a�h��@��z�:�����Ӫ�oa`��X�)�X�j�'����lfď���.�f�X��@�b�9�o�YN��׀+��R����Us��>Cox�|e����ò�i��ܒ�|�ko�]
��.�9ÿ0:^�z�,�?�+�7��cވqg�0Z�(4�`�K������7��}�1���c9��C(�4��S!�3��p���w���$�O�V�oe�E�O�w}�iOt���Go��5'!+Z7�O4�����O��ܶ\!;�}&@��ź��$ś2<�g$m8��O�4E|A[ ������1��a\I/�6�/OvɠM
�]����vY��_��rG-��m1��FIJ�l��0.�-`BxUҔ``��r	�u�jMŬ!��j �W/F��,��*`gq	�r��/^!.L�a�y�e�EY�x����"�'���=���켁�$�OOYf�T	]K�yN��W�ʺ`"P����� ���m(o7��;-4pF��؄�~��r�h܈��n&��beM��1]�|y�<m��@�&+-��5wu��b��t�����zTbM�^xN�Y��v�c��W����{�4���Y�S��\��q����� "T�ϒ�3#t�e�˓P�ܼm�fΥO��^s������扉*�m���>|X��Ŷ�����l$-9W򦉐����l,Q����Z��c>�&�CĜ�p�kb\��x��D�CXGٯ.r�O�J���g��d0=��m���c�	1�^�?�L�)�=⁤�����i1�dF�U����A�����L&!�����G���O��~��@����{Ztm����J��s���M����B)����ƕ����*�u�݋���$�k���GSg��R�C��61����!����O&�%��x,����yG(��;�?(be�w�A8h��Yo�˩QT��l��;��C��NFw�Q|���@^rM�7��Nb
:TA\������X�
ZM�CBoKE�"�[�gN�w{��˚��``
y����ˠ�&}����k2�pa��pBX���`��g�:�pz�[���x���0*�w��轫]�p9IIN�G`,v$ðF�$Pl��"���Y��,�������}�7��D�HѐN�(ߨ������S,Y�99�J��R�1�;kc�y�c��#��ʛ���:_�s����6��
�^p�a��Q���gp�0?c�W8��'xs�PBzFL�Kbλ �jKb�U�몍P/T�R�]���K����e@�k�ə�Q�\%Z'o�����^Y����:6B�k����[kZ�pW3�3<��@1 hM���Jp���9�g=�� �Q`GGő;�j'���!��n�Mt\�	7 ��Z"�Q����*p����03�lW������!?}k�0XXc�l"
��zN��z�u}�����u]���K��<��ci���]�/9��0Le��J��&8�ù��H��t�+Wr�4��[�	�&��B�{
|s�����ߥ"�:M����(���(J��w�c�2C�j��c�A��`��<A�����N�YI��1��QW��W��7��j���>0��Ő��/�fP��ź��w�1��-��u���B�♏���B�"�,D�؀j����pB8*�g���h.�b���
Ԛ�ȭ�������@���I;�G����yD{�ï�2�8g�W�=H~��=d6|��k�({;�+��@Ga�����:������Q��g����dk�Bj���6�HQT`���Tj�)[T���B�L���L.����� �M�9�����bW�WQ���������QEYX��6��9��o�*�ݬ4�A���p�������������x1�eE�͍ت�J�u��؝�� a��8oj)����oZ;��
��K6I��w�/(׃�YI�J����8dI�A7p��k���oi,�j�:�&�h���G����D���@:��g�G���Á���E�z�c�o�{�B��V���lFnf�F����EA�x|�O��KB��b���]gx����\��vLW%�:���k��uQf�$��V%��2T:�q��%SʔS��Kԋ4���rj[bo�y�����Ya�/3�ĳ]^oX5�.3 �q�.�	$�9�턪t��PnǬ	 tT �(�1��C�AL����ߒg3�h�7�3��0��&��*b�*(�#��^��0��{�F��u��e<��e�|�ద(�~ٜ�����6��#g�U|$ܴPT��6�u�a���sײ�5�2��!�7Z���ϕymQuz��7|U|�K ��"ɋ����P�Y��{�b��K�yW�V	 ^�;B����u�Ƨ�_�'�{�����?����|h���vѬ�c��� �"��!��Q��H֘hw
�>=烓��X� mͰ�o����5d���W\X�5��<p�g�/'"�<�3�$��ɖ
�a}�6p��X�����<����c"W�`���х��Y.�o��ɽ�����Gw��	e+K��x�g�M-���@����K#qK9q8���A���� �tc@�Dj� ����I��W8����=O�� ZrOʐ,�ˑϖ�+̵�EOd�C�Rf���;"����_8?���q?�CJ#Ҽ@`+ױ�)A�۠6� Ip�/m������_P����B�%�ߤ��c��[=���ZEN��	�l�hj��f��	��Qܖ�&$��ٰ/���"0�?�� ��(ⴗ"Fk�������p
,��+��8hQӕl�N�R��MR]�
�;zi��49������*�栄{����[��Y�qC� vW6�p���F����D�ϽM�#��K�Q!#�����>M?�F8o�g���(dL߫�?��6�{NON��+G��vm%Z��x\*��Թ�"\��.�B����'¬��e�C��� �[:���x����.��|QR�����Ҿ�Ȉ\�<
�wsH%cOc���:�z���L&�N�Bg[U-��eƈ�[w��`��Q3���G��ZV�6Ё�� �x�bڜb֢����9`sY���u$���&��(��p��;���+�d�.��D�}`�?ː}�@ea�y����(s