��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V��v�8�fO-�6�`��z>�so�B�P��O��W`��^��}��:��g麆9�ɣi��^��(�Q�e�LB��ϷW��ۿ�c`i�5�`��QY�u��$��V)����v�Rx,4�YY>�}��q�L�+u&���Id��4��b�phH���Pr KSpxG��=~���m]H��h�D��b1\X�%���D�����kG,�#4�w@.�tHrx�8��X�}-IE�b��k`����2�!&̡��
��NB����ٖ�0V^c[����k�	�	T����?��*^*�gY�i�m�����y�^���N+�
��8_�T3�� �&��sh��N���PO򅌅[/	 ���C���M�*/�=���S��}<UL����!�q����o�k�6/�Οj:�R�ʲ�tr�zr���B�?����w�m/��]ĩn9�$R�Dx( H\�N�/�I؜+ LSOZ�I��g�!?�0��/��i^�|~�z�C+����5����9�@��*��>@�b�CHzk����Y�d�уB�&0/ � �){^�F8�$@�<����G���K1��	��o��އl����L�1g�n�2�Ýi]�SjI�$A�mCSf�bM�e�[M�4U^);�~��&j�l����EA%3ݷ�_!AaӶp�?�36j;XAܞ&��+䰜)����\���wK�L�d���r����Z���-���-���v�&0|�lq����s�NzR���Nvr��h+�*�Qj���O���煑j�"���#[�ן����l	~+���y+c$X��|Q�pg�@/�oU-|�H�3�D)�co��-(C2۔�T��v�ڤ�	13��X����h�blg��K��zP����3���E���TmV�R��)W�����k���I)O����_M?.��e�ہ�og4���Q}33(��'Y�&p�;�kf�KHiƊ��HM�d�A��o�>�(��<Y������:�n�Y
Ҍiy��82sFU%�H�_,;��ɏ�����Ԛ��q��ۋ,�us��	#��>͇;W����M/�#-@��G$��X�	`����2�N���H�c�x���ʥ�Jz��� O[-F&+�cS^��v}���ρzP�͏����]�cB�[������Aъ|7��LMAs���F�������H�kAI���.R��$������~{Uȴ�1Lߙ���8Y/�n�dN�pN�N����;s44)Vozw�.�C
c��Y��h��)�B�Y�R�B��p�e�MQ�x��R��5������?�+��Me���y�̇]s���Mt���F��m�M�(�B���|LPE��&7��/�fuy(�֍%�ng�U����(���{WUFPs��d��1hh�*�$�;�ᅢz�ꯖ���=�}h�S�����Sb=����ȃ��(��Ye��{����O��6'Q!�o��)S�T�ζ'G.�4:�n�0��y��n|D���;�� g�zP�I��d[���r�-��3����?8�Z(O�tT�Q�Se�D�d��Ic�Tҭ���v�E�����Ϳ���������Р��6���T0m�9�Ӽ�m�=��,�����x�ڰ�+ӾdP5�3�RF�O��B��ݨ�������&�_��s���>����)Rt�p�{
��G��
�C�����)��,pU���+uj�C�h�*��n	� ��B��F�}H�zV�,xm	T��v���If��9KT�I�*�1Q����6b��Nr5<�rC�۸�#b7|�E���2�;�����LM��{�<��]�7���gb�3����y˸��\ce�ɤ��T:�$|�Mne������~X���!,�m��bᯙ<�2�ߵ��*&}��K�JJ��I�X�b�/�뙲U����&e�V��K<d}�OuT�
�ΑQ�O��+|��.�l"D;���}5e�0�>���������qf���M�a٨Jfc�]���qqa;vT ����X&���*I�d����W\�)3*���#��
���e�y&Mw	3P����f'�l�W3��=*�I���3�y��:��ȕ%���3K�u��v� �8�)	g���|d�/c�`���4�l��Զ��o�%�-IįC/��E#��^\���y�T��g+Ø�P�N���2����T0D�?�9��x�H֏���I�p�*qP��R������ 7�(��,�
MJ��mҬ�e~�/�8.R5AMn������FZ�F5�{��x2'At5#�c\X�lb!��BwUeI7>A�jꈫ!Z�G�m��i��L�
�ݻ�+�o���T�4��mͻ�ӎ�ͳ�	��!?!���m�et��kM�����5u�,A�S�E�:U#x�>	��%r���Z��"Y�����<Q
�sw�#�7��������72��x�5\-;�i�~�Ӿ@�%�_k;��v��mX��{T�#j#��k�x�Nu;�'q����E��!��*D�e����f;�0�CBX�{O����R����ˑu֓���X:g��В`�ġ�_����D�r��5������K�e78Ž���y�͝Q�w/�4p���A������ӯp�iqgl�vx�ᣯ<u �4��;j��e��Ptzk���H��g�=+�U�����wAhe�h�U�o,�d��u��&B���pg�gCx)�Pog����hj΋dwd[Ͽ��]�9\���J�<}�>�).�<XF<+]1a�'M�K9\��z��v�6�88�d�n \��������c}�_�