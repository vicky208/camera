��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:�Q�z�n2�H�U��θȊ����w/����`��������pS]~��Y��h�����$���l a���r��"��Ը�+��D�� �ؒ��@�&Z��e;YC�����z�)MT�F.���Z�d]�I�!���7p`��%����ԭ[�~�d�,+�9싕IA��H�~~����DV��ESNp)���#j���4��kS�0��$;��d^Ж����H�ڪ�T�Qv��#PM��oV���O�s�/,�gs4^gT��OuXs��O23� Ҧ��IcZ��`�����l]�ċG�inţ6��4��k��f���sl��r)Ybl��U�I�_y��ODEi��>>����ˊ��}n����g��nܻ��x��Y���m�|��ȑ���Mw
�d�m�Rx�N����ꁁ�.�M��K���^�6iKԳ3�0Y��!��j9x��Ü�;)~�LQm�t��&�3p�z�XY4�r��
�t���_�`�O�G	�ڟLc�B/��rR}:�w[<�މ.lz�.	���)3�f���4�����6�ʞ�\j��lv"��mKQ��RX�xc�UnE�3���XI��h��0����!!��&�z��#_&}�������o�Dx9��f��*��p$��v}:��D��:��.A#�%[�!�F=L�ԗ)���ѭ��������~�������/ 'ND{e>�2�V?�(��<�<�-˭sТT�i��{I��� ʅyN� ����G��i?#�	iEu���B2x���Yƾ����"u�A��H -C�^�[OZ�@�4�2�Bo��=�]�J�
z:2�h��T��*_�<�� �y[s85���g��Y-���MG�$���er�����
���������:�ӥ�>F#=��iȌf�-�M(et�{�DFG��;�V� ^e�M�}�Hp������R8��A�*:�.W W��7�H�|tTA�	��>Cq��w��J�Q�a���&_��i�=��+q\J^L'O��~��>lKH/(Q8haN���0qp.\�I,�<�2��H��1��Sq��ěnZ�Ch%-��m;	�K�Q�y���������ǃq����	u��r�>jSq�Q�o�X~|$˂�ERi�3�BV�1	<z�<��>|߸g8������(�f�pO�5E۝}$6�M��uޑ�^���Ì�@�x���=G��朴]���2�� ����c��+�]��_�k+��o��)���@?9y�w�o� Mt��mF��s��\�)'K�`S�5�=����/?�^��h �w�I���8r�B�,�R%x���)�܂ht�L8> ��������$�k^��)!R!=lO����+p����Ɍ���}l��`� ���Y�s�_�;j�!�}�mN�����[Ma����*�䋣�{�,�D��b�}�Zk��������i �]�[�3Cx!�J�Ӭ���5������(X~��{fd�gpR��C#�;��Bw�7	�n.T7`��f��GҌ�� r���1e��L=�-L,�N�4���Qw��K�t ��H߯�≐%8,&;UY2�)���I٤&�����5C����g�B8����Χ��u���w�053���Ŭ�b��	�D��y��5{L�$Q4��d�N�twٹ��FgI��BlG�B�V@F��t�[6�M6����(`���֗�5�%��_�$���S��pM*i�#aUPW��S�hu|_?437��ō�L3HZ= m�,b�2� �G�*bdJ�`���v�/6nIh��o���:&�Q��ak��Q��[�f+��lBCQ��������G���<�Q��P�Ƃ��E̞k�ǵ|5�X��.Ҝ����WioϨ@��MS�2Ȧ�)�q=}�{&�9�YG}��ʐp�p&���R{7fX�z�#`���1�Q.��� �Z9d�l�խ�"�ث��9����Ⱥ���|��zn�ʢ1�uG�IZ��������Ν"�Yt�B]q�O��ó9����åȸ=V��}Ȟ|%���@�,���%u� ��-a�/�c���lzB\�x�p�;'3�)1��̧p�Z��w���z+�>lR~�K���aRZ~��f�D%oI�^h�gv��h}KmC�0��{����܊�c˧^?nd�$�xYx� ���(>��*�̶! ����kr�=�&π[�@���O5۽���\Pu�)��T��KuE�DC'O{���KE;��F�"߫�2���s�״L�Xޯ�OT<$��jo��m-�gm@�~$����=�Z0ʲ��|���!Pl,S�]����КB�FPnlJ��4��A;�zQ@���t<������%d�����Q��1G��6O��Wg������O!=\���Z4cU�.� �{�Z� 
]�=ڿ���#�+�t�����H����A~ک�������0Մ� �2�ż��Qyf������Xwlw;@��vZ�V9*+�^�e�@�Pcvv�����9����e���Z�WL��f!.L�t��;�"�@��,r��k��Sx�TLcz}U�a�5ؖ��H����5���^y�̤u���
p]���H��Wm)�Y.��v��o�M��(���m�a˭�O�7���?s��A��lx�[cd���Ʋ3>�9Q���q,��1�O�4(��23D�J�󤇑Ж�q����*%�B
 �5�m����ɫ*�s���V��ٻ��R�FmQy_mD�R��]v���Mo�ګ)%�j�����4�1kp-����70�y��85�8/FE'&�yBp��e)���.R��ݹ�ya�G��V��!.���B�3Ӏ���A���Np'�f6mРO��(0�_4��G�*W:S�gbZd�!i1�k�JzT���\!K������8�<-�^�h��=�0�'2��:��|�d�?}��d!�� �Z+S�L� z'�*�t�A��j�V��
^�Z#N�j��[�	VH����!�0���?,�Q%��w2����:�r�������}n���b�O�&����/ZZ�Q���
+��"�K�h�~Z�U�������䦾p'��fU'%%�"�U���ϧ��~ ���@�N'������U���*(Ĉ�bR�@Z�b�F�%c�ՠi<���(�}�#���5ZT*�|^��Hf���k<���rj�^8c��Q�w����T0���#8I�b�=5G� �m���M�:�7,8�i�٧ �5-�b�����ƽ��	��F+���%Gi�&,(��;�=��}�Rj x�l%�~��+�����G �J��5X7�q����2%~8�1w�z�"�%T���d����U�J�|�Ƌhj�
٫��ݏ>8d��< ��@t��p�C5L:��:!$�ǂ^�����<c����	i�Q����Gy�_Fo�z2Y)���g�%.;����e�0�D�5�g#]=~���B�AF��Ճv���B�L'�b�����JJF�Y���V�Ꝩ<�����YaQ1�'8����zt��O�F�\zn��s�@������<�Ս�Aj��~�E�+�x ЛG�|����O"~�P`����N�A�Axg�JV�=��hr4�
�'�E��(+�?�h۵Xv����V3�E����&��qdW"dlO@	,�O-����Az�	�ڳ��" �,�Ԥ�LH��G�VQP���}�d����OOǀ?��"��?U��o�VZ�,[�VDo�v�I%�R'4���A�O���t�a�]�]?��;����aP^z,�jÎ�W��;���'��?�E��C�׺���*��	=�Î�!�΃�A�sSU��/2_N���L>�?6'�H�UkcmW�d}*��a�,C�R�t&@�(���.h3_��`���P����f>�%>`�������ȥ���,���[����T(9�e��"���fN=<M�}�P2�6�B��ոB�f�6�V�"z�#mV�����u�|�ѓ�k9�؆��sm,��8�,���Z��D=�g�ѳ�U׆�?V�#����Ͻs|������&!�!��5�[=� f�-��7��diA�wt|$���ȎF����b��%G�
K����ʺn}C��� Ԫ`��-�N�`��^|+cQ�x8^K��k(���4����sW�ɥ�S�ײ��r{7E� �K>���BR�m�]o�]!˷pt/������ ��r\��*@�A|�s���V
o�j�oB�����Kaހ^ u�U��h�����&qI��J�يR�TO�)�f}b�m_1�*I�P�E&�6��A E'3�R�a�����Z�5\V�/���b��p�2�C�"%��79�ӕ�<A���?T��%p�E��$r��qٲ�B7�.�"� =M�7)J�T������-Ɇ�F����T.�ۭJ8b����I?��cF��4���|{ZW�^#�a��nb�h3bEE��(�N�f��Ct!��EI/c��50����[,d��"�=�{�`�Y����I8���HUн>��M��D�����m(?$1~xuoM�G��4���������!�a�X��>�{�`�$��[��K��WW#���>�7H��񥞵#(���b�p�
f����ފ��������w�yU�ǳ7NO�QQ�$��%�u.�А�G=XL�%U��	څ��;��#Es�6�LX&�#y��|+��_���y�KcQ�l�z�bz[����k�UE��.���o���	^��(,�x��Ё��	�#��i^]�JH������;J ��R	�.�oE�S08vG�-lj@�=Z#� �'զ��0��:}7�X�T5F��tUW�c�����/������+X�f�e���x��u��>�����4�V4��C�H���{��v��>#�Z"��74*�[�ש�9 ץ*">|�}�(00N�	�� ���|ߵ9����t�cqv�1�Q�<?%׵ʐ���/�k��X���38C��d)�/�َ�5�wr�8��ĹYw�$�T�{ �ДY���z�|���fB��2aSi/i�����T�����)ɠ/�F��7�5�J^ٝ!ᷡvЪ��Dd�8��?��� a$���G��`G˟����;
��Z��P_�gz��l���Q�,�ټ��8�ʸ��n���fu��T+%���~�>ɺ��F}r-I�9�['��!v�WB��.8Z~3�d*�Ԛ��O��|�&�ؒ�w!�HܰL��x�Z2�j�K!���O���K�>s�G
�E��Z�
�iI�V�h� 0���^@+�O�|���v�s�wC���%�ҡ�����^�n�6
��ǃ���G���G��c"R��d��!��ѹU��
VF�l��o����ejټ��������\<�ٻ ���C��D�����m����g��It~,4�	N��������h��Z`)}b��sBqx�ճO���K��t��jf���f�=��;�-����f'�tC���p���@�th�X��
�Q���z�7ߒ�,&�!��pEY"F���	�w��qj�(�K "_����←��}C����R|Ԙ채���I-�6L�P�����Qw��z>9�{������QP:f�W.Z��g,��(D��.\�]�I
uE��9�Z6��JZ'=B�+{�	��.��Y��#�������EC��M�Y���A���Ɗ�������30ey���>6X�\���5��}���:��Q��s���J&p���-�7U`���f�0�x�Ṁir���: WAd�T�^gu���n��P]
���^	�Al`���v4�4�Ni�qP�̓�㓼fs�"4�>���X=�3-	hZ�`����0p<��{��#�Ts������/�1�Y��d��4�DN,��2�o4��GQ<#������ZӾ�0�S�d�4��Ơg��.�&��?VU��z��F�o>���Z%}�.��,*��8,vBI/˅��$�IF@��X&a
d'h���c>�Y:��\!$�>�7f)� �UU�ڪ,o���UU��>���3\�y<k�kl"O]*T1�Ր�6���� gyk�qB7�����xgLc�m����~7h�Iā�^y�{��Or������x#���w?���
���]$Y��2Я��7"	��3�Xo��6@nf�S������ |��ֶ����*\��x�dT�F��O%����,���T`�մ&~��ubb�߬('��R@���2S'�V�:�����6�B�o+t׾�K�rT
?O^��>oe�",��0`yoQ8&ܩ��B���t����3-�E72�2�pez˙�����5sc~6{��Q�� �+� ���3��Ey�˒
�����"����g��i�Q�pfE!����&(���B<�ݗM@��x��G�fQ�3�'|�*</ҏ"�ѣ4��]�Z�Fhn'"��e}��Q@�cԿ�3�Cy�)���՗�T�����-ELӹ��X|���@u�}�1VP�U�.�����EjH2���0�C���ٮ
��$��Kq� r߲n����_��\�E5��@����HP=^�
Rn���M�΄(�RO����KH�q��mF���{1���qu*��<�DN���1	g�����W�	Х/��$ςV��mtF�h��L�>�T�	���u�y�^��
������L �N����e�t#����$8b1�i՗^�u���#���M�'_i?�Q
���_�(h\K�`Mh�w
�����h��dmR�ΡF7El<���p!y}�/(�R(a/�{Ї�U��tw�71�z�_~��7�LW�	<pf@k�:�4���o�"۸�wİг�,�� Gk>=��]�ѐ�%nM�����	t�d�F�I��9}n�*C�%�Q�o~�b>~�-�7D��)��,%�	"}j)�,.�=���}:���8���	�ZD.��!��I?��MM:�k��R# 1@�ρem0|�kZa��Ċ|��� �Zu���^���c:W��:0#�Cӕ�J�C��_A�-c�_�93�1X�ٙ����Mg<pk �����P��R
��LG�FEQ��w6����\5��Q��{���'�#\�>�Za0j�J~�+��4R��f�u���43��_����_i^d5�e2~����t$���Q�_��*^#����Ԥ��zX�7�!����V�5$t�~B�8�S}��o[Q�rǞ�i�ѣ%��[`��� �{/��+}b����<>�WC�iLi$^���*���@H�@�{�v9�z	���(N;�&{)L���ő(�JSo��Y�PG��k%�[��B�4}�,�S9�8�X\���#�Z�jP�bPG+��	���wKx�Ɨo����w3mIUZ��y��>��¼�;�K;�$� �:��Cf�SSp���	�#�\�dj��.�#�>ߢ��x4}R�������RJJ�%�n$ޝ4�{�!�8��K {j�?u+�6�L����#M��~�ư��Ow�l0_��0`1N<o32_�CpL����}��G�43ЈT���q��E~�����w�M1����L�I��	�����M{����������b�Τ1E����n�Ǒ۝��Q#���r~��(�ce�R���N�er�D�.n{h@E5�*���'�s).@C��/��� ��Cj��������:�R��^��૥�-ĊU�ʚ�"FFk[N3���F�@��ɵA��j��~,~)�~#Ac3�Dz	��
�	n!�!̡�[�Q	J����o�X�v/6/�'l�+���j���Q�[�V��3★�K��8��7 ��!h���|<
u���t��Fj.`�;h�a�{�`-�7k�+����0���9C߂P�ǉ�~x�D����⮶
�J�<̮��[��`�D���I@V\��L�Ë^Im�-F�6�l�J�a��ޘ�!�߭�<S��t�kE��)7#^&�5������t��Sx�J1�koW�@�C�-�Q�C����y$��$�뙁�H�c��ơ�P�	�d+k�T�&���GP���a|t4)�l�t�;�3ɜY��� �s�r�D^ĳ`���~�(�ؖ[<��܃�㈡������u���N����N��#�ܬE��Y��#�R��=�w����!˺�X�����|6
��+�x|�}:h����ro�'/����)m�aes)���E!��46ou�u�|�� �)�=]}>�5ӾS�w�k��|���A���}B^�R�Z�>�5�ME_F:�N�5޳�Ƽ`�ji54��nj�^z��� �X,;�����2	V�'�7��:���}�"� Q�V��r�*{���^�u�V%)��ӡ'��q`t�XO1���,
�|m��"�$��L+��������T��>�g�-ԑ�g�W�Ә����B�$R"�<$�Kp��U>XU�r��-��CL��"�uv�΃�Ǎ��+dț�APw&���妓.?��!�c_h����>"˒�������K�haF��FaMRɨhm���3���p1�:�i������PX��σ�L|q�C�-����Y�O�e�^+e �8����$�a9s�3o��H��e�HJzfg#��<���JX}M�B
Ǧ�\�^;��܈TP�|P7�>�t]ධ˂[��u8a\'}% |��=[����+J���svqZK֕LEco��]#% J@)AA���*���[[L�h`�nU���>#��]�Й��������IDdN�!�r!h���s�9X�����-��!��.d��#e����A9jA��kTS��˻���T�7��S��ص	�-�HͧT��_�芔Q��pĦ�&Ɩ�kV��������pئ+��Xl�!O�خc9	� R����X��kPDFh��Ռ3��s/�؟�w��"�C�����I{���uj~�bUm�O�e<D��ё]�0Q����FY��4Al>���̊S&."$��	��.v�����WʞdN�P_A���Ҧ�o��b�{�i?�6���D���.�Nm<c�����!��1�nX?�
��.u���;|z�B,/����d- ��7�SZ?����/�t4@�����t%�6m��g��M_:��-z�gBe"tʽ9Kg
�z?�H����>�2?Oۡ�Ea=��dbh.���6�p�����!N�Cv��qV�/�Sd�2K�(��ك$���d��i�m�%y�.C�U�hx�������<�fD0A��}���6^v�m�PE�$�\�lCydk�y9k� �w�.��U[!y;��UA �߀��*G̮��QNBL��:��V�����t`�a�{�۠������: sR-E���$U^���}���f6�Ig@�=�lb�Q�L��=7��˃幬���#��}�9�82��OgCS�"��S�_2t�#�iR�_������S��zA�K�7A�cJU2�`Yڏ����f�P��D]���[�m��3�})7.F����߂
!��@�?s����������Ek�ν�~�	F���m[j.�4���>�D�U��[�!�rr�����O��HI�Ī*ծⴳ�'���	�v�ܱ�����k�QqFy��(�ci}.8���Hm�򌞔�����$a���י���m;8�<�<^]#\�`�!����G{��T�����D����q��
� �����ž������Ӆ�Z�$@���(0�� ��i���))�q��� ��E�).��1>�N��C�u�������Hb�O5䨧�nIy�.ZO曈���l����k3�V[����k �:~� ��ۄOKN��.���boR�ob���Z�$���N�-O@U�[笣�x�O~Nz�1������yvn��fN�5��ږ�Ux��߅��t&�=��G�(�$��L��&B�&��T�p�7BI�����Cm���'����>?�̖/�?H jA�<97Off
��Y9���>%`��Ԇ�6M$����7��me	b�q]��R�/Hj��`�$@7~��p|�V�Ql_Xh:����Ƽ;��b-Vע�K�Jtw�9�a��m�,'=o9�o̜%o�1H�m�?��t���F����ECJO��9��۾B���N�H���@V�X7I2x5*1�C�P��?��s�6�L�O���l��ʚ� `ˑgk6[�D�̈;P�������P8�O���]~Op�[!/��Y�@W)F7��r�69�z@�߆�,	�qKf*P�U��Ǵ�*"��u�+��z�(�y�7iD�?v�9����*{��$r}lU����$����3f�Hwq���]��z1uU�I�=��Űrg]��a��;_�q��Ͻ�+a��=�/�ް�]	�ҧ�BK(��?{�Ư�}��%�e��y]��8��NÉ�=�������{�'�D��PY��=�V��C�9c�� �������a$n�r��al>k���Г�ͱ��8ڏSH����~;ӠW��2�=7�g�K7��W�LA�a���X��, J)����rp�%�Q}8RXu���]�Md}���sŘ�6���XD�rqA(���Qt���(|����Vyy�k�f���M�� 8s���<(�ܪ�z�im�$���WlH�m� }�x��'�R!��o{(����6B�aD������֛�L��9��H%�U���wnI�R���:�ڽ|T.���I���葤m��e*ظn��NG��l����@:���t�!]KD��K�(�K�н$��C���-¸�	&w�UM�v|M�kN���&��TC�P��L@q�h��Ǖ\c�6ʞ�vI-���F�ʐ�I�_�v��⨭�aש>d'������&��Md�{�6��I���h�B�`�Ȕ�Zw[X]�]6�X�����ʅM�Qoo����j�Õ�\b.���"p-�;�`�3x��D���R���=��s-�g�VNoa�{`i�%G{��&�X���)��@!��>X_$o�\�F�k\:�c����s��?>	hG�W��lh;d�ӛ����]���9Ҙ=��i��	z���R�
%Q�K�I�D�֧�]��^z�3Š�O��?Y�ϣ\q0�x9J�I�ܶ+��V��lO�#�&aez��.ͫC8�;�E�ť���$��\��E
���֬����L*�C�0vAtj^��Λ�餸��mU�P��C;�"���0�s�7�
�yWʜ2V�=�΃b�Q�B'��a����>hB�8�"�J�l�Q�[��kw�A�Z.���DU_�ca�ZE�:SD���x"���<�6��e��;�����`5-����� ɜ�U�G��XGa�a'F��
.��[گ8l�M���9���1��,\�*
���2�-p��J�a�~����*4��,Hb_}ਫϏӢY\jx�j��/ެ�RWO�n��Qy�M9d��3$�Η��׉o)�K����W^@��T���2�*s�]`�0�f?�)���ܚW�������z�ӳ6�Z|ԣ��>�dBa6P���v�0fE0:�c�(���P��-	�f�M�Br��]st����e{5� ���	o@�i�r����Y5����B�[�BiZΫ��Mj!�Ѐ�h	YI�O;��A`��A���l���%C��$����W��JX���&�Tm%�b
'�!�'J�:۞��c��6��x�ކ���W6�T�/���Bn�e'm������F�ԃ�+�@2&��!��m�B�W?�)��qv�ꁔ���2Ql8��<�ɱ����a$�f;o�z�|���Ɣfh�Y��6"/�ʍc�6��
̫ڈ���U���MΦ`3�A�V4��S�H��_~i�J�N�)����v:�����߯�[�F�ɧ�i>�۞��bG��E(��y���:2+C��X���)A �ա�y/����)��;�-���Ky�]�}����C.{��L��Z?�D =����,R��!�
�e�߽n����v�z��nt=�w��^��A�:<���Ĵ�I�%��v��ze�q���<�g	��t����� !b��$��_�U)�/$Q�E=�j�!+}��O�S�Sڲ67�a1��o�uڵ����%����[�K����\�å^jz��t�KˁJ3I-a �H�:���ʒ؇:�r�G��Q;����i���#CNN�Z����킫u��?e�z��i���2��՛�px=b����	�Љh#���T*�.[_Q�L��?�p�RE���7Ĕ?j��T,5Kt-���3��U��}�@{BI(����
��;)�,��gd�g4������!�Zt7I,����&O�%R��2g�md�V��n��Kh<r�㡊���<��U%�D+v�(������QJ*�mմCgU���V��1	.�|���u�j�%���ո�hI#���Vy�C�[�����uE����"����V�9��B��N��M�����^�J�h�傄��) B(����Oy��_!�89�o��Ι(O��� ���/��e�������g���@SBB
�?��\�mJ��8�ˏ�"��Z(zٓEK�#��\���M4pc��n�3d�wS�Z���jI������|@O�Ѵ֯6�f��s��A�~����I����@s���x���`���� D^0�%�[.W�AI)뭉=n:�˗�E|ϯ�g�*mO�
i�x&�w��m���n�-�������"����n1;U`��3>����O�{�V�u��e�cfQ������=��.�|�������C����@�в�c��Qr�A�b��8�I)�	�0�*]&t�1��p4��Ѝn��W"�
`uj�r�O�lw�~�|�vV,�ꤝ6�V�K#�U�$��)��(٩�e��i� �+h�;K�z�5&����Dh�^�[뮌m����g��!l�����aIb�Ƚ(���?���2~y����|���#D����mcH+1�p�·^��OS%86Д����Z5�-B{U^��5�'������ g�gxҏ��=8�v٦��t'�F � dE�Y���W��H,2�"��������x�M����qs�ج��?�=�H�pr��7�Q�"�,��hgy0��0{P��O�[nc.5�������7q���ap�P�!�q��)�ɥ�5]/�w�������3c���т)�	�+�����9�A�:K�0��	B�fŶ�yo�m���T�Jc
�R��U��o#ʠ<5G�#6��)�?	��!*�r��e����i�O:�%2e���ř;RMM�8�/4C������vr;ƶ������8��^������B�>�>J�ԁ)���3|T(�dώŬ�w�]�>�ה)NK眻���2��+h�%\8�k!�f����.�֚I\������4�!�������k'_�Pzߙ>�!��O�]S�b�Q5H%E���no���e������@smS9h��M����y.�����2�P�2v���k��mld�A���>tA�א�[[0t]��2>�o&ӄ �(�� 5	��L*�>���Gx3@��t$	ɮI`̓d:�fa8���
�Z�6a%p4*B���´�^����,�@j��0m9�Hy���j
�� �C�ȴI�Q
";X�☳-X}�'��OA�M-�q���/��:�Eۄ�k�X85^�}"c:�h��9���GW��5e3U�
7.}�|�R�.h��n�^)�\X��)]DYǜ�Wؽ]�70}������a����]\�<�]
6Q�8�
n�k���KJ���P���	E�Ez�n���&(�P��8{��G�]P�q���.9�<���ύ���P�m��'<+����V��hK B�C!�~F���������ܿ�;�@NjId|��ՄR��wM͆u������&7�#?L�\��Fg7LX� ,�s�]C\4��;��>�1�aC#fvE� �C��u�G��o-�|�H&3�?�3Z�>�|����`���@���?Oe�hx	��]���h�Γ�D�H��,�I��mɗ��99����LC�S�c�.�c���g-ǌ��b�=�V����z��;���٨es�$�D��^�$�@#�v�w����Bg��i2{7��ʹ�ZNeO:��z�C7ِ�g�~��a��� |��Ϙ!H�����$��Tu��T�[,Tʥ��r��>;���>˓A`�þ*���[-�n�BsV��Ǻ�bXmAq 
���&��lm���hXn�Vϧ�bj=��d;} �p�0I	�d6���wsq�j��PR�=��z��o�<o����e�?���^Wp�}��_'U�a�@�S��H�����g5{�6{��rh\����8*��|^[ǡ�?����D���#�<ޒz�r��տ��a��*�;���_s��/�z6뒮Q#�*p�^ޞl����e��P�rn�[v��*������u�ɤ�4�P;�[Ȏ�aY�)y�dWu]`Y>?��m��g�Q�;�����ٙ!Xِ{�o1�
O�U'�o������R`RLW�DQMx���� �`�Uϣ�+[Ņf ��w�+�.eDfF ff�(�E�r&^u�I�$�ĻM;F&��c��������T��{�T�[kl�ƣ�֕D"<K9^\Z��O�!x��~mV
��
Ɋ贁<�R�N��g�:An �l���[#IIgk-��%sC�8qj�/�~�H8@_^/���5�����5�
Q*�1��� Й<~���A),�kR�uÃ�L{;����=!M}�?�/�������u�>u7�5��AU��}���p��쟴�����4�f;ٙ�Y^�_.3˺�"����c}�A���ݽ_"}ѱ��}N�n�u�������3Hu�� �T�ƾh!ܭ']���-���I$����Q����]���*y�+p��U�u���c�d���8�B�E��8�f��ӴY*bΈ��nf��^n$t��c��(�dWs��ܩ�%
7c���"���|�:���'���l��
���t��~�lF�¨�t�_�
�^���7��%^X��P���h�f��P8�{u�|��q�`ؙ��/�14{�m_�JC�,��f��V^Y ����y �ޓ���&宑_��Yg�*&5�����o��|�<�����(��V���Y '�z��f�E���5c��юRJ}h�������u7/�9#�`r�BIN�<\�����E�eP���hm8 :�9����H�Z'29���1l]T.\���F-  h.�+�eEH�Q��P�}�M�,�9�q����m���J�Rp�#:�5�_V�CU�
�}�76��:�I�^��`T�q�{)L�����m�	D��g<S�.�^��{��tL-|���s4T�p�����^c�s.Ɓ�O�p�6�� �)6tvJ(,�,����F�����'w�]N^{�x����	��4��5� <R7�~pp3�I̟h �V>����|މ5���s��r���a���@�# �!�T�K|`���[b�5�-x-}E�VE�7�&ģ?BDnP�M��ly�%t�k�c��Z�I�qVS��l�Ӟ�0�Y�:H�����L=[J  �B�3ņ�'��ف{�hDo/Vɱb����fo �̓KN�XVmMZw��WGEZ[_ {�Rm2<�w�?�R����K<醱�o/�m<_�Qf&,��G�j� UQ����4Y���#ؓ0'"W�_�&�%~lv��r?'?�[s7�;J�t���j���qBT�q`I\e\�(H�d��Ƿ~Y7G��:,
��S��\$' 74}RF,��I�-��Ҍ �k��]�c�+O-J�RK�����*b,��)��/��h}���q�Z��0���a���Ր����}�@�Ϙ�Mw|���w�(�\���nlR{
��g��澻e�SG�pz�Þg�n/	؞�`2ſ�������3�ܭ��G4���Dʪ[�ŪL�צ�;�1��.�`����$b7��;� ��B^���H �����N|3���ꕴc���U;#jo�"��)�l�X�;��(k�OX���=F���%�����x��'?��hr�W.���>���g{ 9Q��}�Ss�߃�VX%��[��T��4:�����u�%"8�d��K<T����Sb��"����Y���@��ఈS(��d��`N ��P(����$�+-Zp��mP��!���|_,9��h1� ��g�������Q$��<<���S^����Z�pX���+�wϣ���.�E5J9�p�˃�~dG��������I���=
&%��[��}�"�9�iKE/H�M��Z�b��	"��!�$\���<���-����H�o�{Inù&���Fg�RU(Ƚ��)	��
F�	�(�����@#B�89�1ޣUD���C�� �b�l�ڰÚ'PG��ߧ�/epÃ�C��Jb�W��G�:Q�)"#��PT61I(�������&�ƘkHWC;�ʲIR��iXP6?':�����̋H����ܼSrk�b=9~��~q�g_u!�2�|z����%׈�+�z�����6�%��W�Qm�\��9x����#G�`����z5�t�i�_��6��D����K�h^�hi���xTX)���M߉P��Ss��i��u��)�� ]b�q#��7��:����4yS�2&���\ߵ����4Q3�-S�9(� Af��}�q�K�I�ٚ�WX�HW�;�F��[�i���3�/{ $�w>�����_tfȏ��O(e�~<Y������)��9��.�o0C����H����-u۷γR���O�Jx���6�⵷��U����,^��]z�w���$e���i!�@ꛄ�3���J��<(�>�w
��abȪ(�*�^���1����ul����ew��vȦ�6�W�ASpm�	���c�*I��]9�o�9��B5�����H����t��\�(OE��%������g���GA�Vlkh�#���G��,���G�β�k���~f]T<��ÆcV�̛���'e�i)xs+7��c�(p�쁱9�pi���]�VH:
?��#��+��Qd2�ї��[��nߒ���S�����M��u3W�QAoX�H�M�I��D'�#��T�����Yݤ�*�} �c����شR�J-�?�Ko�W�]��rQ\?�ʀ�	�����pMnSzQg�G�p����!X�_���c�P�>(J���=���)ɟ�v�V�h��_P�^�R�>�!Iǧ T�iq�M&{:᰿�ySP_�%,C@�e(������:0��.��6����d�i8%��0��[���Zp��c�g����h����ܮ��r~�z��YM�~ѽST{�P��qPm����y�5�̱��Ȍsͱs�g���l�� *�M����B��#�T�9���/�>���3I!��Ot�����,��	���Q����s�!���_��kb�:�H_(�X�	��B)�^�eE�^��}1*t�r���~ϴQ�{`p�Y��O�:b�$	Q�Yp�w|���+K�a�k�I���O�Pb\�ܷ�^&>1��8��7��W'O�%���8�rf\J�&:�3���2�rdD{+t���4I�`o^���w��#���f'y#�����e�Vd�JY0��x��~%f�o��3�B�R�%�o͙݇��e�{�Eb�@�z�rj"51�X|�Y���7���!�� ��7�r��� y�hU��!+0�ZA.�971R��D!�d��>����7Lh�K�����y�M�#;&(�t9�J�&dÌ>N�\IM��1��`�֋D�E�ɧnPr���}�mR1l#��6�$И�Id�/L��p���5�Lj���Z<��GGʣK%.��o2��T�؆�
�K|`cG�@��Mz�S�IC
 a4'5H#�R����N��z'1�}�.{X��߹��`� �6�ÓO0��
�G
86�ھnxs�Ip+�1�	�LI�6�[�[*vY5 CȽ��w�c���+ZZR�%�̸Ek�O+��2!r^`/���[�|#8Ԇe��m��j::т"���ޣIs�ߜr�r�j��,�,צ6NVJT�����wK�bA�3y � ��+�J-G)��}|����Up����#�i2� �LDƞ�7&��O�8��u�:�zϳ��S��v����!N���-졭0m(q��Uj�҆����r�-�y�=<~��`za[:J�c��!��s�b�Av�)���`
�0�=3��/��:��4e	�f��IĈLῶ>�A糣�#��v����_���xeA!J������^X,�^P�f��j���3�]5p��^��x�i�J��� +At�T�AJ/��3P��(���{�7��f���kZ��Q��ٟ��(��F�G �L�;7�o,�6��{�� ~4�	fo���D��Oy������l���!,��USC���.���� "�ex�t��f�ۋv�<�%���j��]���Z9db)eGz9�m��^<Ћ�I2b��=�4LZ�����0֒��T�Z\Ì����ٕ�|������Ie5lV�^��������g�v)��U��6���[Q,F�[��
�'��F���ydY �1&���{�!-�3H;2���_}��
T���]�|��B�!�H�_�b�w�����������^��l6���Y�&0�*���`�Laq\�M��b�`5G�Xd5��H��mD�I�~���(xj�����a��=-�;�k0�j��n�*>�y`����5�V:"�̻[�&�M�#C%�_؄��Q�M��f�v��(�$H^-sx��A7Q���/�T7�<>�N�_�EyY��R�;��+��q�����踿_P����L���!�j}w|/	��n������q�l�W��9$�?��~��s4���:��L���$�̨6JΦ� ������VW�hA K���'�{���T�jt���2�i"��!�g��"W�=5�������~�C� }��Bp�;�Lf�Q�6@�Șآ>�6nɫ��g�U^FX����r�~�
�ev{g��9�5��?�e�
�����<
`z+�9U�X�:��N���� �;��F���[5U׫BׂN��ճU@�}:�_d��(Ds+�N�C����4����Q�t>��=����b[��ٹ+���Ҧ�i\�$�m�m-�-�i��P���%���թ�X������x#8{/­�W�$� xrs��kAN��L�d1�f?���K`W��-�|YZ��o*��yL$]��4�5
��>�.5;��$m�T�[|�ł��8vݳ'��o��x��-�vוAސ�w� �Rʱ��g�k�IƠ7�lˠ�Q�V���i{��F�g����k����/���1J!,�J���Y�U¡��~I ?�F: ��`~��F�`l��4+�!����IH���>��5�Px��aJ,��ZuA_d_{�67��� fj�������Ѭ�ڳ9WM*�	5yU+��3��/��� L��ҳ�8�r!���X�B3�!7�J���3^�
�@��NeOD�������k���>�ª7�Lu�U��x�-��<ͫ�?��\n8�DPT�a-�{Q��1�{d4�hs<h����UD�\�6�L�B鯔�l\0.9�ɅV~��4�8�j�e̮D7�(��=l�v��B�,�7㴨��1n�/��HCr���s���(n��d�ޭ��S��kEa���7*��	p�YB�1������\���8��@UU��l]��e|���]s˽�*TU	�t�6q�I��ճbD�5���V�j)������c�zS��ދ�kXH�B �Y�Wn���~��`�?y�֤�m�>)����8tsZ�-9�+���V�+�h:Yї&֗XvP��w��3/:�ځ\r��ٞ�r��{PC����Z��Ir�<�f.B`	[�xQ}tP��~#���W'QK=�A'�; 7��S�OH5{�����
��Wa ��aY�a�h��p�q"q��d}[��57�l;�gT�0�����1����n��CJQ�Rف�j�P�v�S��1����KPVz���T ��M��e�O�iU�����J���($S�h���vg�T�O��!R쳔����{2�����{�C1�K�%m���F����������Pn�5Mi8��/�b./%�~�i*��@�掲���nA:�sXʠ�hCp��,���a����[~e1ϸB���qGU��z��Y��2�.���[7;��X���.�$oG��/o�Kۯ1��	���L�{u�Y{�W�cT�A�<M>��c����w��C� �3ȏ?��<���>���� K*h��ɿ�#?��ʟ�/f��Y���0�Z^�fb3��l��*E�ׅ��L�/�c�
�8>*+8�0~²�R4J��԰��j?+��V�y�kRe�e�'*����[NCr�"����[0�2R�I�z#A9�/\V$-�N2A��ev�'��qC�N��ۭp�ٖ�ʖK;�Ϋ�k��w�x$=�z+���KBV�dy�o� n ª\׼�YiQ@�f�9"�̃Du6��ǻ�$��@��-n/�g��eh~�%O���Y���'�{��1p�5�ʖ�"}��,�vh��$��OO��*��hDAbڟGPz� !�KZ]Yo���Z@m�W���G����D3���U��u?�����_��������Оt�u���:�x��~�md��J;�;�E�T��݉4��~�S���4Uc��4/)�J�4e�)a΍I-����|b����{k�����F�`�Y�x*9���X���YO��D�r�=�Cj��s��r���Q���D��RZR{�4����L
gPsG�n�h�+_AJ�I��Xp�Ǐs��=�
�wP��G�-i�3��+�R�ɴ��m���l�c��~�݈41Hs�JcM���#�r�m��KV�S�*�ؼ�	Έ�Y��n`�0[$|IT��D�pǈݵ�f�쓢�k�+t8����@��D����{d2��%��4յC�+�A��Bh]��9���&��ɢ:��	��fJٗ������J���Г<+ro&�F��hX���)(��'`��S*u��BV���!��PĤw]�V����!�PGe��?��J,� '�{�gfm���- �t�*N��TV_Q:�Y��}rΝ~� N����\�������W��\�a�֨5ѓ�<
�L-�b�D�þ���9��a�%z��$��IXh̕2"�r���\d��z�!8�%U����U	���K��cup��lF�Ii�MQ��_�6i�Hcd:�^V�P�HQ	0I����O������ Of�� %P��+�=f?�V�,��067wwY� ll|\��Zɒ_�FIs��d�bd�B.�G�N�_Yv�޿h}BZJ(�����~w�?I���\�1�h@2kQ����c,%.Zxxz@�!ט�1m~��{Tn��詝/�'���4樰TR��xO�:�`�����@?G�z�f����:B�y�׊t4�W�����3�1������2h��d��$h!Y#!�;>�	 s�8�M�F�Z��˼��L� ˘�#@���H�x[�_�ߐR����aĦY�gt0�䮾�)z ����*6ז )~J�=��>����2�`#3
��!�=��f7�~2��J�by���rn�/S/�s ���Gq$xu�����Jݢ[�Ȇd$e�y�G�i"�h�Z��p�0P[V9��lQ����=�a�_�}4��`���/���@�`d���q!�Ì}�V0s��]�Ej��e\����B6�G���k1�Fhu/B���!��l��)8ݹ!��28�y\f�u^�|�*	3���7>�qOa|ɵ���W�m;x�>�}���#����]R3̴��n�wҌ��犠�+~H�D)��0p�z���_^�!B�����hAR�o�!)��e*a��YS��o��X���KMr%'Q=ke.P�t���YQ�p�4���Y8�sۓ�
Yr�e���<QP6��;��_@ɦXT���)�%�o�,��M�+4�P=XH)p��%�j�,��|ɕG=!/��]�]�(�3I�
FS0x�/��/ѳ��d�K��9�麢��(�>��
=�	G���!u��;qMA��q���)b�r�����3�j皪�A)���b���C�=B�.���B�{J�.F��=��7g �`'�G��9���93�D�S�"22=��X��Z)}Mu��`���Z�.��}��� ��J[	3QW�=�W�=��?��.-o�h�߄�"	r�E_�0�4W��L$F�I���%^m���w���pl�@��X7��[xb�*;�&й	���M���z��Q�sȻX#	X�W�a��]X,��:��f���Dי!�:�;_���}�O�|0��Oy�q�m:�s��5�~\��5"&�m��o�}C%2`i�sw"\�C�պƏ���*�g�=E)J�1:��|rg�đ7èbh���9G$�P�K�L���`zK�Δiom�N$&U[ �Y�\�,�_��}��io�����!'FA�<B=X�|���$rC�wV�"��u1�fƚ+2�^T����r��'��`�z�m�OA<v�i�[>��]΂�<6X��G��Gr��c��	M�;-�L������{Cg̔��I��s�_������!��J1ؽ'q�<� ���V��@�Bh��ʪR6H֧$C@�{E�W5�>
���	��������k�1���u8uߏ��u�I��ʖ������ds�NX���j�C�7�d�4طS$��c�ݽ�����3�[�ȰF� �������}�&�!E� �	IQc�!�����0����[45� p��'���5?O��z�E�(e����o�+đJ^�$�7;����PߛM�H� Z`i���`�X$��N����^Ӏ�S9*��7`E4�����u<�An���"���T�i&)QE���킠�o��jK��n�p�Ξٹ���'/�{�M"!�� ֵ�g)v�׬x'86���ݿN���R�	�5�I���'K����R�g�?*���N5scT٧.�郡����5$B�� *�\Mn1-��6!���C2f�L�����c�]��P{�op���1C�0`�j��_��S;, �<��F�$���{�/����䠧[�����aT*�:��(+���?M/ƱX
��r��K��J��D(/�@Ux�����$��B	
ۡ��{����� Pn��*x,%�
]4?'�0���6���D���g�p$�v��{�s3�� 7�'5M�D��e�w��6)������;u �Xη9ޔ�m;��*�C��K����������
�\Q3�"4�����]x�Fڝ���+W���_�{5d�wnB�+�~6�Ꚕp��6�5>�a��q6П����"J�o���S���Vĝ��Y�"�����9%XX8��0�x�x,G�и�my5f%�s/l�b�xs(�I0�P>���RX��<8�A��k�w,�k���4��:{�Z\�gc&����%1=fn����f5�/�Rn�=�NZ��@Hْ�;�8*����3��t3�y�E�4h�Φ���@Dg��̥��@�?U�t�kF��C�D:5 ���&T2r��1��\f/�)��$��
Ы��|V���45@#
�B���c	�H�LE�?�-���1$c�������P�!�C��x)���p1"�Yu{�ˏ���?2��y@���F�7��oO���>%oho���e�F���(���A� a.`�s�'8{xo���U��v���ʜ����P�@匰�\[��~̝��E�VAsH��u����YW�"6'@�6H���R��v�#������D�ʄ�ͫ�����>����K��+ߗl	��wO��-���d'o+�A�h��q���6F/�O���`�󶭱@�P=�)]6�\���"$<�qmW]���I���*R�	�40�M܏h<�-�^ƺ)�����k���U�㫢�A��w�ze�g��H�"���g�H,<"�X���hG��d�E�G%o��� ��7��qc��ײ_B�*Lt��#h��l>�w5K\�K�OPAo4C�i�HU�J���b���(a|p�9��k<�o !7�&̏�y��k�u��%?k9b�ژʖ��u�5y-�e_F�~������H�͡_����c��<���3�IfôD2߭����-8�c�;|~ػ㗓�Ho�i���^4͈G�I��v"�K�f6�O�.����9𣫎X��|[W���s8�}�A%�ƇoY��$g]	��RP����)��[ <�hl�3��=�W�U����0��BLƀ��e	\��͡�g�c|8��B[0	2A�Q��+ǒ�2��N�����e�:��w�Ȣ�8���7�iyƲ�+Y�����:�}[�&�0�~�t�M��Q��1��#�ՠԛO�X�|����i*߻S�7��#�z4���JS|2;B��IBO$��sZ�9�Z�4_-��-���ʰĘ� t�b%�9��C���Hj�;�~Y��ʽ q�Ң`Yi����H�7�t^�0��:�R[%�L��O�P����pѡ��w���� ��Zf�揀��=����h�̯�����ƁD��Ǳ�qw�@�B�		��nR��3��t#N���0��rЪ�M�x���Y¶��(<^� �-������G����<(fH?k�%_�a�o�`ٜ��˸'�=�����|���#yMK&��(��s#��KE��z'� Ȩk��HY����+�Q�V푪 �ͦ����㝊������Sț2k�`0�Z�\ 
�X�}��"A�:Z�p!�	0�4,)���|q�@ S����C ��/ѣ  ��i4���@s��8>$��{xcJ����A]���~���V���|��n�|�b���������8Ԥku�� ��l���^�T�J'�Ẩb0�pOt\�����[[�� !9�1��j���2����e�N,u�ҿ��/�*��b|��"���.�� �äS�B��/3��?V��m$/�m��p��#��� �C�R�� Q�X�=�
�(Z�T�тn~U9��ke���3����+��<"J2��sL� ݉I�^GT�鈀���01��MU���8H]�X�&�`Yv�IK��S8.������1�r�h��N1�@���w �~W
T�[cg(�f�=(":���TD���`��z�S���]��yل��r���97�<��e�"�4eI��x������o����+1cîp8�_�8j�dj�&e�R�$��GWň/9%8�q-t ���>M���T},�����-P�Aυ���1�Ow���S�|�]��ߨ����wJiv�̏�� P^#����=/U8J�Ƅ_'J�&P��b�#�>+U�q�$��9ج,�j����dZw�d��.a��7��X7��Yl�L�Mt=�������y(�Q������hAq�&E��U5�8�����;|��g������G��|���D�8�0�'㞖�^��^sL��qع�#��Ցl�=��Z�	`�6�����ׂ9�EE�A��.�xt�C��ޖ#��F����M �i�e��i%"�m3�$kM�]Gu�|$��<��j�+�W t
{ J�mf��e��d+-d��R[Ќ�A���<��Y�Y�s���Iާ��u������8���+��rz�@]�};�p��Ӫ!����w���T��d�\�r�%Q!���>H����35]pKc�x�wľ�B:d,������2Ig�Qu@��0�d����s��O�@&�v��>���$Rޜ�&��jWKo4D���\�"^�ȇ8�y۬�R��9*��"i��假���ԹJ�Z�j}��yN�2Xδ��� D
���3�Y?� �W�
(�_�va[��%\�yR�	wQ���k�3���r��4c��$�jmÉK�֑\)���IeDcv���KF�������k͛�J�M���R= qZ� ������?-�z<'�H��"�33�Wq��F8Xh�������X�����C�C=�з����y��⣫�g��ȷߡ�LO�_H�&� |�*������c�e'hZG�9��7<�w��Q�g���V͙�,��a����p����I�\bC����!�Y������t%��r���������brV��vMC,���yʃ��A%���[�n��r��gvx{i�ׯ@NL��w��Ð���A�e�)plw1�B�xL0Fm���4c"�.��IJ���_%3��(OH\p��W�|S��zqp��$I��޻S�	�)<��?�RhS�m�}n��Nkz^����t�+�J�'�Z��铸�k�RR��c?/]*;�d��hƫJ�S�D�G7V�|U��(�^5�S
/M
f�|�N�j[~�]�7�ؽ���}ǷphE�)���+�NN�#+A9��+a�ً�1nl^{�$�}N��ƞ�)��G�@����%�"2�K>��H3m�R����!�^H���,{�İ��F$�v�(¡&G�:e��z�ꕙ��*�ҝ��d�G�����7ҾE�j&D�|����ᓞ�'��>	��x�u);��!�u��A^S�J�+e}��6I*: C:T$x3ڡ��\��"d &��k|���֌��i�^��oHb�''��-�oW$C���&H`�ڄ��>�)��(��ƃ~U�́5کúK�+n�Y;C��1�SH�~"?������g�����(��~en�P��fb�׆_iH'&�ᓖٮ�K}����$���p��U<`��AǊ7�}�/:�i�O#�0������+䩔0u�,co��l�?��$���:A�g$oT>m�������!ZI���>����Ҿ�u��L��A$�D���̇KU��=�Þԇ���C@�P���|T5w�;Ye�8Z����tG����I8��¢l�oj��B�?��d"��k1s����\R*F�i�{'B�d<�j�"T���~*�.Y�˖T���E���E]��(V�e�0��[@<�k��KX��̸8�,Eo{��[���d˥� xi�.,XB���)4��, �wg'�$�2n�������c�c	���@@����F��@ N�W����Gc���o#J�v���	�̻��+�(r+x.U�����`(Q���V2�n����s ��aB�B�{�*���7��*j�}H���#"�j#���$��L��XU�r�_@-)�YF��TR����4�=#�d���3n�ƚ�>A�N4�Z��E�DBH=�;xlD'[��)��w�b��I㽝*0��G��J%>,C7KڍB,?�����\��y���t��]�b��� �mN{�a �۰@�boވXt�����<��l��0���>#b�Lĸ:��q�r�G^�[0E��J�^��rxޅ�BL{f4�y2���FeE	ר���@ɷx �M��K�������'�Z�h&͙����h+t�Ch{>Y�9��sa� R7�����=?����IC���2d��]��<�F()���yE2�1A�Ȍ���3>��H8���8��
V'��Oؓ"ٕ臫�K��i6��+��,�i��ӂ�d�ez��0x����Ҫ��b�о�Tnr�䩾�`�C�x��d0�����lVԥ��|<�; �$�څNK�$�V�Q=�,)qu?�1w}ޥK�`P��9U���R�X���?����o��Y�d�^1N	~��p�^CV��tO�.a�������g�>2�_�Ԅ�nK2�9#[�D�a�6��?Ӫd"�%G�H�_e+���e��|Ѱ�9��>GJ��Ҏ"�����vʫ����Pf7'AreC��� 4��a7�9}��h�6����_�y�P��\@�y�/��L�gi��\��]⩩w��S6�/�hٵe�F�;%�E�O)[�<�z����bTlJ�ӟ�z⡘��C��$�q!��jݯϹ�$����V�yl��z�,�{j!\�Q�](�3وs����ap��Cf�_"s��TEN��j��ig�K7��rS�����Z!��E��X9����� E�N��B�����Qb���ߢ�5*�.�x�?+4T[���A�5}�f[嘯ǽ݉[��P�g��tS��7����?=*����U��U	z�^�g
b�7���7/V���~iQD"[�4��6z�ʄp�y/����:�<��L.���	B���s�ҿ�Z�@��8����M|�E�+7���;��e8ʥ�Y�����+Z&��v�;Hx(�w=E�@ۊ陞6�sj$�i�o�On�/�R`��t#?�h�"
����mv����M�6�R�{�!K�w2S�Q����;#	6�^�l'�Y�'n(~���	Ʈ��C�Ah_*��}
��a9�I&ס 7�"��Wi&tv&��rF��lΣ<�Dא�����������X���Ŧ7����#��OIS��)�JT���c�$T��N��4���d� p7��Л��{�-��� �t��'�ÏM�x&aw�����"��
�((�;� ��?�_��	��Peh[�6&h ���Cb�@mT�]
�2��i%���:WF�o�(��i�*w'���ߤL.,Y��0ԕn������Q��y%�ғ}����Ζk��ȩ�K��Y��v6Ca�?p1�+�a�?�j�OvW���Uz�'(��"*:`
ET�-�\n="�����|��j�|����G���)���A�~���C.��=�ռ��@��'�۪&���^�u����m�-G�镁��Y9��pыj��['�o�z�y)2��;�"Z.k��	l[=f�,{��h�NZ9��T�9�A0�L���M�@�3r�*C�-�͵@F�10}I��ef��&�~v�D��wG5��+L���������qA+;,�A�t���,�	��칬++x>긜YEYz��� y��4>(5�-C�����4)	bO��cx���%�I�TrOO��{U�Ai���8��Dr�`��D1�:(0k�b"ђ"�DǯC2'����`�)�N�˗e�L���W�R�۞╼GA�Gr�;֒įa�a�)j�i�]K�	� �o���J�DMD��Q+M�������JVA��pb��Y-�kѓ�^�0x��as�.�)zcWn�]g`�a�e��%u�f�dqUa��O�h����m��{���V�8���ą
Y�,�f��˝K�>���<�^x6�]Y���6;���3d�T��M����)=a�[}�	r�y�����KY�o���-�G'���d���~h�`�ȧ��0w1Z��%qkע�Wm��Ϻw��
fy�_Ďg�*bܯ��*��pG1��K7��cC*�Z"�����d�I��M����L'"�	)�a)�O<����_�]�Ж�L�ܕ� ��@`����Q���0*	�?�n�<+�aw%c�HN�n��Gk=�T��a��fٻK���e��'�M��o���d<*��cÔ��<����xk�t2a�Q�?�G��얎����:���K�t�XP���0 �fw�VB�_d9'�!{cm �������4��
�N��e��P�\TH�>l8$�>�B9�/��<���pR�qd&�F�f�E$y��Bӳu�P^���PVδs%q�6/d`��)�d������n��k�b�� �ϕ�q���S�tϝ}b4��K�]4~��f�	�}��Q�=�}�P��N�����fWzڣB��%&�Fry�]~u�4\u|Fڢ;C�'�/願b*E���
N�Z�SiE�N�K�2Yz���'o{�Ƶ`��5�A/n�����w>�����H�]��+$���X�_���;>��3#1�	����=��\ZNz�H#��@A�LgqW����%1K_�3���cn�{�
��U�)�U��J�C�"*���u8�M�>�Շj�3,.��J��y���) ��5�[�IMJ�����^�&����v�U$���.�QS��uz>E��eo��@�����!�L����c�sx���|��.3l�Fpq���C����ѹ5�����FΡ�|�s'�~��O���8]��Q��cE 8�	ߠV������
��c�G��o��<t���Z���3�i��Ђ ��v�݆]�HI��f��L �?H�u�_g�۸~U�Z�vY��'�+�\�ao�D�@�`��鹱�J����j^mϑ"YB=F����N�b�ln�p��c�-�=����C}���'ɕ�ٞ�֪,����&�2��$����ZI��"*��`y������kF�d�`,<l�&�J!��յ8�j��(Ĥ$��*1��̋�-i�O� -�o}~���z4���пt8X`;���S�6A[��
��%hV�j�f'2����s�_�F}f��'~�����E�Wz#|�ύe���R>���'�l�ה��7b�fSV�a�uw�V��F���F�V� 8HT�Z%�|}��;�1�s�	������Y�j�AI��.I��+�3�!�2&����Ie\�Uv4��_�X�#�y�z`��D[쌌�G�����|�a��yö��u��a���H��Q��a�}9��a��F����W��������p߾���'�L���݂� ˴w����LJҳVb6�u�)�a��������#����u�Y�[��v���A�a��^`���_���+o��[��j|]:�'a���l��)�Z�7���9a/g�:�j�����2��M��	'n�r#T옝M�Y�Hp�����NsG���q�7��� �g�?rֹֻw�8��$ �#fvL��q��I����Np��9!7��Z�Xt�!���2%T�γFҥ��g ����_���<��x�!���EU����Hb��,�)mi1�/=(��=	��=&�T��%��UAķ����ܠ��x ]geMI��n�e}~H�0�����kÏ_u����S2{98(���oh�S��
*��^ґ�ҝ���T�]Z�A�<F'�fa)
�_C,��_��މ���⟹	&��Qs��B~���,g�m_���y��f�W�[o�#�����lb�;_��n>e�I���9�%��V�AP&�+3�"ID� }N��ih�<(�S!5:�$����3��j�ٿ�MY��T/i��o9���R0��<o�s件�'/+0�Sopff��	��3���Ex�q�/������>�`��Tf���4�?�L�Q��$/���y��K11~b~��8IIS�r��Q���0�3`q?�E��mZ&fs�D��I&cE8q�Q�`��E�q�w���C�},� H3�י�Y���þW�cb�jDnK��V5��
��@����"�#W��l���	}+g�(>�D�)�Q�a��Tv�5��E��_YC�����gYQfM�a6S�A@;��/���Nd�uރ�Ǉv�d\跻*!�Pg�>�I{BySJ�ۓ�㧣
�N�^�\i�-��-57VT��5T��5l��y��?�/of�]"�˖�y�G� �n�΁Y�ݑrZ�B]�k"P��@	��<�(E�{ȐW��y!�p�����U�EƷ^+��W}��Ws��U�c�$XK�p���%�<Y��Բp�%/�r�F�B�Y��+ē�fܖ�f�Ց޳l3�4�A|����tܟF�Z����dC�/v���E<�l��D=�����V�J
��aWd"�0�a)tV���qU)8�L,�L93CƼ���{��A�N$� J�Ca�ȲZ�2#<��m)��Q�6ΎVfx��y�e��~���I�_������\��`����|��fН�-����aAO�P�������Fd�;��Z�)&B�LO΢q�R:��z�����e���,��*��Ukk?���h.�_HXnM��3���BQm�a�����?Y0���ğZ���'�8�Qs�t�7��լdj��jh5��s`����7r[~0�S�R)���^8o���V�� ��_�_���Z��(�s�.�@Y���@ntR��U-eOl�>�O�!���b�	./|��uCO��3�<% �y�,���*���Y�R�t�t&� }��B5�}��!獝�!Gu)�8�����/�|y(β�20pr]3Wm�g��C$~U-�~L�������a�u��Tg��vh�~>ɟj��_gh׌Y�=�^��o���g��)����&o�P$:�Y6z�F.�U����,��	A�� #j��I|�� ��ME�W��$�+Ȃ+�ɝm�S��v
'��	uX��<iokw\v2�ɺ��L��7��E���͜5sh�\�$�8�D��}�Lx�
e��9����j1�QE��(��v̘bB)p! �4&��˦=���g��静��;I�.���l�����;N���~ <A{fЀT;ͫ��; 7*�WR�if'��.ʁ�~|���3�qԮo�r��x�%hn�n�@��#R�N�5����=� �	H���NJ�Mi�
d"j������n����/���X��י��ǝ.h��)j B���(�#�CO1��G�2^�TJh��H���Q��>rs��IT�ñ�.�О��[~�u�i����>�����Y/A(�k�' �S��O	dE�oI��N)\^��D�ŀ�$��|;]���=��u��@U� �qs��\�J%��g�G�1M2<����I�E5�27��j�BT'/E�X�T�E24����h~�2�J�y+x���ҧ���� ���Ğ˳�F4:�����Ly��'z�0'Z\��Yʃ�륂q�b��!�����4���ٙ��&���9����{�	���,J������
:���tX�F�*$\^T)�=\���~��^ŝ�%q�k���n�lŦ��$+����I�?R�����MQ�W1M>d-_����,�����{Ӣ)o���|�=0�~K:�aaa�R�+��LSs�Z��2�QQ���_����O<�Lט�u���s���g�Qs��.��5:1g��0sZ�[ѻ���ٯ:�dI�|���a������;*�u1���4��a�sl�}B�ą,�#����xC������s�K���2��^��gg����`�lq���Q8����x�{����I��+М�d�o�<L+8-f�h4��S�χ�s��?am'x��|�s�3 Be�@+Ձ���2
�t:����r�X�<�����ӵ�y��Ȼ�BTvU�0.5bE��{sfP�ߩ���[r5
�$�$.���^G(�u80�1���)�Y����2�����	i��M>oe-&�� ��� �M��^2C�XB�Э�h��w������|[d
�lk�k��8ӕ�v`��I*�4���Q��9h��a������+��j_�{�]/hs��C��vGBJM��$�_�$\c�A~ډ-w�}���l1P��b����qgK���(Y֬���(n$E{9������iSګfH��	��gR�D*�o��� ��p�I���l�ƿ������~���Juc�O�_b~.��4Oc���9��x���v����p��d?��-�CP�$`�r�/��#.���Fv�֕�:/i�Z�3h�d��
�M�5?\�$�����kX,ڱ���Ќ]�[���ĢȂc$�z��#OL#��	�>}��!
%�W$\K��55�(qERrA=���X���{�������v��D����.n��U�x��3T��^�H�Hu�����F'oq�żz�=icr �P�5ϠT-�m�H��P�G�?�+�\�ѥ��Z���F����e���r�Ҕ� 4c>^���I~.�Ct�e�"k��q�ۂ�����}Yy��r����H���ɣU���G/�I���6�%\H���]D29�1��])ϳ�����@���c��P��� F0,{:B�uOfq�+D�����7>͗��o��N�D<zi}G����W��w/�ά7���*�g>��[#B���Mۈ)%�2ؾ�zI-��h��֋vS���yk�R��D�iSp�5���$�PCi�]������$�>�LC�7g�$�.^�cw�38��}Bu���F�2�������jOAv��eWQp�:i$��54�4�U'|�'�DY��$�M0ŅG��&"��Xo�e�\_�������x��"�*�������7�Ղ$98�f��@Oϕ<��T1��9AƉ�j����$�c�[)�9�*��U�F�<�L�\!�
�����ʩZwKa�1��& �r�\���䑼t?����)�#'}�
�^�ln��F�7�e۲(�HW�X������y&�<�	�&2���0��f�>"�: �~�#$qã*e&��G�Ɓ
0x���B��lro֔�蓬z��^�#�B��
���M�y��=�;.���=�`�*^v���Q6�VɈڝ��`���L�����!�Y���FBòtGٕ�bi�����9P���p�@,o�Ԑ5�bX�w�̤w9X�g������|�����I�=@֫9[�N �iվ��;hOp1�������g�c�ɘvӦ��L b<[��Eg��&�+ �>�!�v�F�)�O��
�>�vqw�0<��tW��O{�$�=Γ��é��K?����hD��8RI�1��3,�s�}f��`G��9��O��f�x�{�ӎ�Q*�5��$�<��^[l��aoT�3H���L(�΢*�ë۞�9�{�!�^F�A�"���b��� 	�FAH�%nU�/�¥�g'���
�\�i��X����D:*�&��N:/��ֱ˿�7e2�{X����ڼ�[���Go
�Zw���AKx{Ĝ�b���F�[�����C+�'h�BA��X���2�k8�-���U�H-U�#����HX�Z:֌h=�ms}���-ja��[�_����jfv׋$[�ɬ�W^�i��[3����g	�P�)��:�~]G��(z(�c�`3��xqeQ�����y�����e�5����3�r����*W&j��pMʝj[0�-U��n�1�z��h���%v������n+���x���[�`g9H�蝎���*ʀњ��ڧ��T��B~��#�~9cۡ�*$�@�>a�B���Ʌ��]̑~���X�&ҁ_������,����hR_�����[3��<�f�7.���5�}jA/zp$J�QAJwGv@��2�
%���B�j����Р�Ay�4*����c�K�L#��v�PR�S*�}�U��d\�`u��&���b�l{*�ܔ�ъ.O�>��?�����'�D����^�0���}<�~�b0���bc�oUt�~�wktq�LK'��?1�#ۑ�Ї���r�{�1���,�˻s."��ҧT������@�#R� �x�#�]*S��l.s',2"���Xn��x�s�3}����Y�.�j
Ts����k9����9@?c�oZ����),)4�q*W�כ�ة�AE�v0D�\�:-=F�B#��pH@X�@���f��R�%q#ё4���aIȐp�]��1C "�
��ͪؠ2n&��o�%�&��g��f�(`�_3��Ѹ�'4��w����[�NK��qj
�煳4;�=gv���|�U*�C��Vk�����0w[���.sJ��O�vvei�+(�����c,A���5�%(�3s� ������u�ܟ̔�_�Cч2�l%>0��4��ʥ�h�~$�RЖ/KH���|1K�vʫWj^�l%)m�Z��q=\��
��zRd7D��.u4�oƁ��p��������έ؞=!� ,w�x0Z�����=NN�h���LN�wH1`���V(���F�8��?��/4N����
x�23��BT��oɹ�����"D)@��*G^�_c�^�b��9d_S"�PɳLݟϪC���ff��޲�W6CA������#P"���?n�o̱O�j��a���m�(�ۜ�x�BƧ;wE���ێ�.W�hF+'v������$��c� �i5������Å��Ǜ�9��[(pαX���5d���/a��t���r�<��B���0:��.��[�y:v��G�O{�~��]�����_�!��}�6�^b���,\4�\�#C����`6�Y7�Lp�b~Z����#�Q��	Cq��X��#��ft�p��q4���r���?I{$�$>�G ȸ~��� ��\1��9��������b���tkzLZp�pᔯ
�.��P�S�Ւ����d���E��"b*�����;�/n�eDU��Ǿ��rEI�u�F=A��g\����te�n�����(6
 84�ܰ�Z��~~�cƲ2���o���	'?^�
��[�;�z��y����c Mj'�k"��О���F�(�2 N�8#clFے7�������䳖�8(iZ�蘫2K����#U�ۏ�P�!��3~�"+�mB{S���e����)�~p��r��˼�M�`^§�ᘓVK���m4�hθ\��L�!L��dH��Q.�X���0,m�$1�_����^l4xdgMu0��LG�ML"����
K�l��
��A�|7��OLܔS6q�c9��sD���B����\Ƨ�`��7� �ȳ�xu���D7����v���\g�;�\~ɳ���pjK�����Q�t�Y���jx����n�fU�7����V��dˏ-�ph=)�fR�ka2W$<Q�L�ξކ�^ź�t�����8rÕ1���3Y�$�ѡ�N����Ʋ%���u��I��3,mQ `%�^��f�RtP���)s5��P/W�j�j~x���%�ʾ7��T7��o�^�����u��Od\�sk\����_Q�[��b7|��F@��?���ZVR��ȉV��P�uS�u��9� *�ی�1�-f�f/>?3�'�Ge��S7a��>�& �'�g.݅���:,�0���jV�r�/����{$  �?	��@Ƴ�P�����U�� �[��$T�YrY&	;mܓ���ƨ�nKi�Y��_l���P.f�М���划������e�Ş�#gu���o�3��)�L��O-��������Ϋ0~�g��>@�GVY6>��&���-�K�9�੆߉�h+�Z	�����bb(2��Ex�I��i���'4 e~Ȇ�@^�Џ��q=w)]���uKm�B̽y҄�IJ���#T�I�����M��[�������o3�$���g���¾��^|��Q�|X��SI��+�ˣ�ߩ��SKN��W��]�y&7�B8؋��q�p���^�F��`m/O��CܷZ�#�n�ZF�Ӛ_����J���_�l?T����{ ثvwT����H�#Q4�S��_��8��vh�#�n���
�5Ȋ2yy'����|�Wf�ًE���N�����LNw�U!�� E�W�⚍Xދ{��ކL#�E�~ZZ�|3iY\�����jc�%"%���7_�NR��psVY�C*g�&K����I��k`El�#����`��;^w��.]�7�:5 �4�¬lFJ4�k&/��]DY�5yw˞��Z5�
:�.��"��f%9*��}N��р)�o���jS��학<��PXV\���!���;�#��d#�љ���H]t@��T���Bd*��k�Hgh��}�U��g1�8���53A˦���M���w�p�'^ǡ�5U� �V�U��nKpYaD��XE���oզ�7j�ՇG9z��F��A�=A'7�B�S'�,A�J1����L�����e/�B�g�ԭ��t�w�/���)�_���0��X�팣��@�@ex����@�	�hr�Q;��u��ԧp����(q��e�s���;�e�<���;
�L�~=�E.3q��;VS�7W��2�u��C2�p��E���d��i�������y;B�͚��y��xxӲIr@��-�� V3���)rwV�=F`
V��ִf]f�_��s�V�.�ǁ/l=���do�	=L[#&�`�r^')�:�.�Th V�#��~=?��?uq�t�����V�L2��:�g���!}�=x)�{�{��1nl����a��o�6�>��I~�j$7P�5����=ԑ�����9���BI*�.�A��*�~4#N}�N�_��)�����6v�>��fe�5fI�I&0G_%R������TO���l�a�Ǎ��!�G����u㭬ϿF�3B�̲��;���1`5�������Bm�����u.�B�Ѝگ��e�|���'�g��g4jQJ���`���:,�N�*O�*K�ژK��ئ�ĵ���'�g���{�y�>�ߚMmڌ[7ݩ����/l��B;��ڭ�&۳�kp�z�R}*:'=��5o&bb>A+�u�����O�~�Z�p�lx��i�G�K$/��P���1	e���G!�T]��K�.о���Edp��D�+\>yM�ˑ����ԇP���{����R���,�������g�I���*qqH�x�	ąw+o�CP�D���\\��wxD�e �9wL��}��'�*-�����B-MSh1�x=��J�L�m%�Tso��F�OX-��"r9����䐣M	++ �m�A��)9�[�x6c���*��կ��h�݅b�O����|��.��)���2FO�s(��<�F�tXP�>� n*��p�?8�
㠪�yPY��܄o\�!��d���Ҧ�޲�4�#����g����Ty�v`҃��d�$ԻM����#lHӦ��Ӻ����'��YL/�Dto��B�?T��eZTZ�`��ӭ����lw��W)����砒��X��|��2Uò���Jlm�/���qČ��SO����{Ԫ�9bW{ErJ�d�5�	M�N��}��4������&ힸ�H���j hx���ONB���j�'���K��K[��-$��gO0�Wh�����!��c�m�E�?��(�{�N�E�\cz��:�V��"�
Aο�gە�j~�����I��8ͯ���$=5gI*<�ޑlzm|B��X���	�%��ݴL�m����pi�|���x��\8F�M/l� �T�vc��]Xl�3�@S5V'���b� �t�;%�������8�OmG�s8���#���L¸cD��?,��֩%A #���8|���!RF��#�]�}ϫ���^H�j�gGI"�
�o����f�n�ri�F�.�����Pޓ����ɺ�����|I�$7!q����bp\ᱡ�T�YRzI��;��$�]E#�:���?H �w��~��3��	�2ڡ�@P���~���y�TqRWAPM�e#���$<�VN�Խ�jz�}����=S�8�W�c4(99��]+�+j�3�rHcG�T�XQl<�ٜV���r��������|��
{�$]���Dq0�Q��uOq���[Y�P��\N3����4d����h���"Y��U>h�0�E��n�S���9�N��M� �+�Z���=��${���w"����ܿ���|��T	��;����?�î��}uwlS����ިN�3�p���`�1��U�F����d���l�K�9S�o���m#B3Ȓ�M)Zy�E���0���O�3��E1�-�us_q�����7�y�(L "�%�¥��p���,���9"i8瓽f0��?����]��E����|"|��%-v��t�Ŀ�u�7O�`��3g�w�
�Y6ढ��V���Ĥ�����Ϲ�1���g�G�T@��/�,��P�E
R�>�GK�\�=�H,X���MY�Ī��M�X���Y�{FRe&'�^|�
^�Ӈ��U�-9�xvAJ���v��I��J?~|�q�����xf�F���g��S�-���@��D��%���+M�+>�h��.�<xLy� וn����ā�?��R�yJ�c�Aq����\sl�g��V��T�?���W�1��9Ղ��bK%�dg7��d�L}73C���c�*B �P�i������n��fαB��ھ�7o\+��@�0<|:-�J��Z�XHHP}9k�becJCuz����+��R�f�����Ij�P=ᖘ�0��?E�8�*d p�I�O�r=-��Ć�
����H?�Y��D1��kùCZ�y�����i�y���P�}-���T�R�����]�������sE�7�*����3�%��4z�GÕ� y����l�����
{=��xH��t���=���2���������S�N��߰�.�C-�[�9!� ��p,��w��B;�"��`�ɥ�bn�:�k8!�d����gݤ�2�DW���>k�X�~��U=�5Οbe�]kW�ˌzF�C�[��~�(�B';ꕔ��!�VRSn��q���֫�嚎�)��Ȉ#ߪ@4��l'u1�Lk��om�r��q����dT�����UR��H�	��=��7�����F�� n����n���ZFHQ1�>�]���*��!l���x��9���y�r���(�Jݘ��Կ�;~�Ǭ�
"�ֻ��V�=h>���)-�s(���tJ��,ףX>�TD6	���Rmۋ�CQ@֤���[�ckfb��1�?2�@�v����3C�Ǐ�Q��yu�s�����/�G�|�����3S�C�-�	�Vn���[@:��h?�x��|�zCK}>�ב��F���S ���<9�圀���3K�]@��E�īVI���͍zb����^���5�w:3z�WsՌ��h}"1�G�>uJ
�!���;SL]e|�7&5���V�\`���^v>D�d"8�^���6�3��-~}��&��ey���׭!��/�{~̂�/��̩".%`6�{�uj7�}��5�4���cH7�8>��C�q���^#d��j3���>�* �_S�:�`����Ui��V�����jG:?!��K�o� �1c��ʓ(d]c�Ɯ44e��_�%�k�)���G�����������|Z�%�-���e��މ)MD��i��<t��X���ԅ���ϚhcWS��h�n�4��(hP�\�f}�1�)W����@yU,��Fg���!��!��l�Y��*ܟ�:��wX>�&$���޳�m�@�_[�RUx�1�ir�0����s�}����tVj��y�Rha�5��U2ӝ��N:������Y~���0k���V�� ��ͪ�om����(vs8�(��ı����S�Xz~�l���������v.'*��Ϩ�辞�tf?oX�p%8w��J#���*W�)%�,�c%���]�L�j<T �@z�����M�s���e�BP�f�p/+�������-���Ʌ&�yr��q�t�/��� ����7�Ѩ�$!�I�]���c���Po�:�n��!,�3��2���E�V��ڈx��5'M����o,���na��Ew�����B�����g����M��,9E�ܼ���f �c��KP�:�}c��X6&�D���ČY���6k�����ї���2�p������*�`vh��x�RK�)^�pM&C|w�'I��l;?xe�h���<@qX��7��H�Z�̬��yO�y�m�G˾�����_!��W�����w�Ӝ��i��Sj;S�L��!��$-)��p���ұ*���o1[�O��ZG�y�����4���*`S)�����k�ӷ�2&f?2n=��|�%�>�Ȗ��DX���z�c�vDh�&#N��a\bs���e]�uw7���_[�|�ݖ>�J_N�רO\�Ymwx��t��q�*��+��z�g%X]��DL�cfs."���>�qKլ��w��7X�P�0�B\ ݬ�R�|�<~�^^#-R�r����f��X�bE����I������9���u��9���Ut?L%�~�^
,N�4�K���L��Y�������GC%:�C�c#�؂%N�'Q�I]٪�eq;$j]@T[c~�X=��-��R���d��R��ϫ���K����`n,tyi�9¬�$����n�AU��:�1�|��=��I�_�-1zҙ���Kč�����l]�Jn����9@��~Y�h�[dtp�F���n�X|�$��]=\����6Q؍��r��糲�|V�}p���_HLN�+�S���V~�-�I�T�Ą���*�Z^b�#T�p�N��mzO�tߩ	.�3�'��Q���q]����w�k�uG;Ybg_Xg�]=G���@UK���� 5��L�BȌ.و�%_�-����Z$Ŝ   ��=�h?3��$}�r��j_n���T�T�Vr�}6	Q@���1������Kw%�]�AL� �f���l�G:)�"��jb�)�H�U�ɴ�}"
�<k�h���&Eh�X��k�`pz�9��R^-�us��bJtP$��z���&���]�"$\�[v���B�����mqR���`��*ܖV���4�4tO��%���#c�r/��j������k��&Yh��C"�B1%Df@����:\�	��=��}��y�\S:^�����ο��@qh�%�e~*n�U�c䴌Ф�Cl	 � Cf�=FU]�$W9�B�-�'���g;0�Q�2��X?�B���`+�>�:4�T�]H:��*���g��3�,�����}�~���k����(�����T��ܪ���~t�ہ�����8��3n$����1���Tf�w�xj�ع�1��|%�'?J���p�c[7�S
�P{����	��FcP�3aV#']g_�D��{D�TK�����!�&}��㐈���"# �-�;w��ڹ�.J�ԃ&\%GzI�x:�]�L�Q��8�Y���3
�g�0~��%���W����)�2)a��g7W����y���d��&�!r`n��ϝ5��"�������d��gt]q�;��Kd�B��b�r��p���v���s���Q:{/� ���6=�����[�W��mH��@V�,Ee������&]�wbj�j=��@�B����T%�n�\\݌�6���ߖH�������P^t�77��0T��B���H��ɨ�k���3��ud���5�P��9����u��P���b�tψ�̭�$�{��N���1�֨���L#..�ri*�R��2ў�dl��*?|Uv�[��W%9������X�����Q���M�T6���P�i$�V㌷�����~�5<�Z���(j�b^�g՝!���d��?%]����=��^�6h���;ߺ}�Qq�q�(Lq���/O*������n&�R����p�'�����xy!!�1p'����s1]1�8*�0ѧ�f!(��'m�5|��pqd��+�Y�������x	oE��Nx�|~���]L5���7.��kF4NIG�M�u�? y�3$�G����}����H�B�Wӽ�-7q���%q�~1*1ll�T�	jS���i�1���N�'軁�r7�ft���D���X@��}Ș �xD#XrҭV_%Y�L7��)cC_pN�w_�Ag��p��` �VwK	w��w%��<�f5��o3l��#{���c����ya��{l�2!�&����L�b���/^�Z��e�q��%F����ڝg��G�i�����[��:sIk�dݯ|���`f��-×��ڛ��I;��4�5V�{ֱM9s�?� %Ě9ɣ.��g�,<�����Mc�8YcF>.���sWu�:h$K�S,GU0%$�ۧ��� ]��u&g�[�d�Q�C�pf6��l5�KI�#��;YCa2�8G�uY	?�E�M�A�>������b(�>wޢ*9�+���i����؍^z��2^)�& ���h�z"з8ⷶ.[��ʴ͊�w����@�sH��C�h�oG0OnO/���-M�)<uܘQ�Yd�V��;7L`0��հ��36:_��>@��DQ7lҷn.�K>b��X�S�<�OQ��	S�Ŭ�=�k6#��_�3� -��MS�{o[ ��ŮJ �U���70��\6�Ml��o5�c�?i��� �Q$����G\]����0��P����|�h8�ƫ
�u����*ᐖ�g���Amc"n>��C���y�\3�*Ç�;�`�N���3�������]�b��YP��'�b��PtʥP7_�� ��.�������'������d��қN�[�U>Iggr��[����0��
�*[^49H:����*p6z�5k�ei^6�M�Zd�, �U8' �%l]�����^�M��wYb��C��kEw}�#l����m���}Lb{	�~�zc�lM�E��R��qV��܍�5v	W�O=��[�l��QѠ�,�Xp-ϥ��T���-�c{$�o( \�?"�Dm�����I�	��I2j���Q��Y��u�ᰯ��mr̀q�i���s��^��8D. �ko�(�
��]��bg�F��{��|�>��@����h��-�� m;=��]�,v�EWA��Γ���_�����%�(��d�C�.�	�r����_ék�����MQIҢ(���f�r�L&7�FZm�}�VT�@��P�;�`�oe�~�H�с�~I*�{���ϛ�	�{�Fc����{	��rs�VŚ�K���Sn|�hDO�̯ہD��j�gx����;~0⅊;����F�ӭ�'8N1 w\Q)��(mo;l�%���s����,\,��a�b�Kv�"?c/���n��'�t!�,�+�;V����v��73����tc�w�7j�u ��s�k��ڹie��A�� 7�����#ײ��N+'{�V�0���;�},�ls��wWl�/�#���S�F{1>h��囯V�αFyF��*��}q�?y�I�4Y*�˥��j+Qbxie>HJɼ�w�����[���B�,�a�h�ZhY�8������Y���)��a:����{H��֐�(�/��-�>����n�N�V=�-�D�sFh�}ߺz�N��Xb�'ye�db���4��h;��4��{\��@/xQ�莵�/����c��:��l��H�x�=�sJn��� �?	��'�d�DOU<�{�Z�J�1��É��V2|�)�><̻�n��>��*�n�an�d�d͋��s�2@���=&�zF����ojۘ��Ə|�;�$c/I�9)�,&;��Q�3�0+׾�ߣ�V��h��T����ȉ�9��}$qƥƤ,��]��O�����<� N��;���	y��K����<�����FJ�HPI*)���͙��u�O!5�Zd�D�`ItD���	�+�`�@�����V|ߠ<����,���a��ϻe.e� �H~����3W����}M�>p<��1�9��|�{����<�ʯ�����4�wB� y+2UM�6�ؙ=�ʰ�y�C+ �a'M��3Fd�I��V^�C��l�[�x���;���z��X�U�r�#/���eet�;�x\�Ԙ{�}�N�`u%���]$��R����bL�R��餍��Rz'Y@Q��XΖ'��[����S�΋×H���Һ��4OF+E��u���1u���פ%/&)�(�R��TP1�6���M�\B>�=5[�yS!���AT�����2���O>Y�8] )#�z�*K��P^d�N_������Gů5�$���P�f���"n\'8�&0
E��}�d�d�&��ў�ip�?���:��oLLU�+4�ǟp���Ë ]���hE�5�>Ͻ�����5��UUQ(����t>3^�;+ͳ��HD�Ʌh3�gz돞z����6��Q��i�OI��\[���<��`�f�Us����1���j��c����P`=-���{����_��8Šl�޷��u-<;۳ea��+t�/�	�Y��>���pٯw���
��u�3�������z6��B��X�W@53"kG��)u�][G�X�f�u�9&3 V��m%��b":����4b}B*�A(�fq� ��)8aٗe?_��	��$�1&�͖]t���tkۜ뷫��LĴ�����]�M�Ʃ�[w_�~!�d�
[�L�q5'G���.���5f�~��AV���[�a���	��l��(z��@��gh���&垁�L�<:�Ё����NƮ/��	�j� ��3,[����%�%�]?�_	
^�������Ep��pi�{0B��(�D힆���o�����d��,a��K'K�}T�/�C��R�|�.��ݹ�E��3��^m�H92�"�
�������އ�&�N6Z�+n콻��r%�j���f5���?� S����RT�7~�D�s3��`�����;ѩt����1W�4/�ʞ��ղ������A`x*�Ƥ��&Ϻ���U��X��1�o;��Ԧ�O�X��$�+�M�e�d�{��n��"�I�{:�k�}�����ۓ<n��=9�};VΧ�]����/�:9�+b\�,	CS��#���i�_��?Ad�Ҷ�_�Q�ǧ{�GV����5m;t���c�!�X��tNC�����˔׌WC��$ț 7��q�*!RN�]�[�S$î���ؑ��Gm�{[(�����d�Vh���-���V>��h�6��ŕF�|����S�y���ьW�Z�چu�1W١b#����/Ր[^Z���dU�^E�k�P��nD�$f�k:�ID�����n��=� fF�<9���w���q��f��Q���$�-���91x)���\�Z�0�8��;ZE��yQ�op��@�{���]C�DK,�X�&V���7bn���#ږ��p���:�K �;zX'�@��P�2gyH"��4@�������Rv+	�6�|�j���;]�)��� �$�A�Y��79.�0���3��u���*%%Iz�S���U��NϹ�_��)3u��rȝC���!��O??��GQIL��L+O����^�(S�[����|�(tN��F�[�Q��?��!�C���	��X����gsCòl�x�R�����b�x�n�g*�&�/UJp��}�A'��@Hc?ܱ�{hk��t>�#q�&+`�=�.�4��0�W���m$���ɪ'����^䘱�7���:��9xh�^<	D]b�'˺�y�5�`���o�϶Bjc��^�3�s��Z���t�
j�d�s}� �ۧF��,D�4���[��jX�xo/8���|����'L��#����2�?̒ȱ�RE�X.�� 	�v���
u������iO�$�� ��s�B��z��ʙ�7FXr�/�1	Ļ3�6�!����qIBeenHz0�qyE�[��V�C��&�ݾ�`'9\��{��V���Q�g1�.���y%� q�|��� ӏ������D�V�/��� ��o_� w��]�d����+DM�a�	��MĲ$D�ջ�lk	}������#0�����p�GlA���:IBOHD�hAR�.$5�>&r�ɳDE�=��Z�E����'`鞎}�[@���Wz�	KC"�9o�zX�	�KҖ!;�|��^��@����s�5hQ��:M�xP�9���,���p�yu$��媫XP3gp�ٳrC����za��=�?��N��s�X�����=��-�X3VE��r6��Y/{�洛e ���m�U���1�N�[C"vRL�p����b��n����SX�Ɗp՞�@h��s��b���Km���l�4�網��ހW(&�����m�Q��İ�mx)A�#/>u>&$GD��@�	
@�~�O���<
4�c�w�rb׺z\>jּ�u^������/�s����M��6��E`���*X�w�:;�PÔ$���*���I=�\���^Qdd��&d�^\��ī`�����^�ee��[���m_��ڑ���<c�=#�Yza٥5 Oֻ��5+�gR�?ynk����x����n��4)��޿1�U��G�9�t��H��:*ck�b����I�J�+ji; r��Aø��Y��7�Y����/2d�Bi�ዏ$Կ����C�Q�p��!ԗ~�:Ǽ,�#��'<�+�P����f��-��k�k�*c���)~�f;Op�Z�f�wwM�E��7	�-��7ze��.�T͸�D��|:K�@�H*�ؕ�ץ]�Bk�'�
�?�@r�3� ��q�iiqah���o��g���3,Z���+|^�8ڽ^��<�e	�SrT�`9��L��="���e��y�I^��G"K���!{�7I����xQb�����	>)UeW{���c�㋊��j_F�� ,��ϡ��<�l?�{7���T&��	��Ӈ��#q��Pv�%�Z>=���sR�����v��R^�����E����(z��C���3����=����xo򖅡�j�p��ب��F�K�i��d�U���;[���٘7b�D}�v��8(�())5����6-���!���V�ފ������E��>�����4��Z�U�y�Ҥ��i%1&hB�)N�щnq�0c�?�K|�8��y�o����w<&�I7D�+���3����>=1*>yP��GbV�@S�7�W�k�O������;Ϭ]�>�`�܄*2״�������W���L!��F^�k۔��;�v8�r�!�+Q�\����Y�2(O�i��F6�UA�Z��~�mз�,w8�F�]���na_��R��#	�o��T�-4B�.	��gE^����iեB����8ۀ��t>���3��X�(���<&�H��v��rS��iNw�G�{ɚ*����Rs�g����	�����Z��f�NA׌!�X	�����&�/H��n^ve�b���õ�]�
�e��
�{.��,&���Sn�"0ճ�j��Vhw�p�ۋ�A&���UC�z��Z>��N�rX���u@��8���ۡ�?7���͒a�&���S>i�f~�&�g^��kv}ϯ0Y�?��L�/��N������h=��kלf�a"q�9,�k��ș��ǃj��z��A�\=���p��W�Lu�����[	<�grq�>2"�U���Q$JnԵKӪ��0�D�>db]��_���
��T
6���6�SO�(�3@�����42��IB���Q,$��L7t�5}L^�����c�g���X������D_ c���YX+�n����6���o��j07��0��2)��}.���9���g �P�H{��C���%�٫A�4N?�/������,��u���^�#���w���JJN"K\�l6u?��8oU�o ��D6��\�T�aF�s;����ܺ
��d�3>�Y�N�I���Nц�ы�.�����I�<�Ζ(���1ܕ}��e��AN ZW9��kw����U����S��A[�F�0 A��=�.��vʽ�IGv��y۝�/�Jwr����M��l=���'N�.�\
�>T�%���F���̈́H�᪠E������~�32��Dovew�%E��]\\�O���^����Y=?؁<��V��{��v���۪d�"t9L� w�\�5B��bk�Wy<p#��7/O*_ $/�����U W�ױ֤C=|��d�\���|ly���B�z�!q�g��Mu�Y�����?n���	2��]�tR�<��Cހ��2���M�/:y�����N�怅2� e>#w���P�W�^2����[�(	V���Ggqq��yz��z���r�����5�U
h�{}�!�S!n�m�JAc�k�o�)�b��?Ф�j��E2���4���2PTn�D!<�ÁE��JOš����}�كT�v1ΦxD���#���3<V��t���Vg��8���/�f���S���Yx�Ef��Y2�>��a1�[��L�AM>����-P汷˘ś��i!�k�:B7O}"��tұ�b����g'Wv[���8�:��cbq��UF�&�g�U H�k��
�p��5�B]�9)���iƼ���w� S�@$�� �
��R)vɨF(yO�Ay<�@���5��;<�6�@� o*/��x<�6��N����΄c����$�^�j);�:�<�
W-R��ũ�t�pm`�@-e�h�rhM�`D�K�,��.�eKkf(�S]��1� ��0(v��o1�f�}׉a��z,`l��ܠ�5Sᤛ������/̇gHI�}l�{�����
��wU-�Փ���n俰�u} -=�k�da�ѝ҅60cI��.�_�����~y�!��1���x��8�.�w�V����N�h�{����ӷ�?��Gs=�w�]�l�j��SP�z�X�fp����q߮�����کC�ԘDIY��{�M�=�4�O�G�?�(�CX�ن=1v���_G�k`o�6ߩlO3� #�w0�J��5��x����<F��&?�X�cp+U���ҙ�6J�
��
�:���w�mN��GJMbco�#����'.2�l���xJ��ZBz���¢��ˊͤt
;�+��t�{EC��[��߉V%��[/�3Uɵ{̗���&�.c�q�>1���^�Ah��-��s��y{�i�j?�,�I�B����l���0��q�o.sIP@�����]�*jc,3�t�Ƃ\��(�8�	�8q=�Fb��<I��[VH����hv|x�C�����u*?8�mq6��c�=�������N��1OʻCI��f��U/[�8_�v��vɕ�k|$c'AV�En�|}�����ČUo�W�	��Usz��j��#̦�6�=�l�j�t���m��{�L�D���%t2/�!(2q��DA��7c�IRj:��~����m3-}]�9�����]2�Z�s���|��_�A�Bf��H�
{62X���b�ogy�Za��i�h%[q���+�/�t<�I>�ի�]5/�c��/ˉ x�/�n�l�g1��q5���Cm�������܀M��8<�|����	���I<���9t���ђ%�:��w�κ-�zX)�?�sq%y%L���4#S�=G�c=T����퇙�2����r��B;�]��q؊�`��7��9�
���l���^SE)���������痙���b��^O l�oD\)�¦}�ʕL�Q[�m�V9Yy���%l���i�������k�I��M��I���uI����[I����n@W�y.��,`�#'��~��{g�&x�Ǳ�Y���R
�q]�	���e�`�{U�z�S�3Z�O�����f��瀒�=K_��Y����g8Ŋ�ǲ�w����t��k̛��O�HI��;[$F�	c3��q=�Z{�YM�j9B��C��%�����Q+�܏���G��̵%�G<s�zM�QǶ�?�d[G���H��Ix�H��eS[�#p���;���v���c�h�H�c)4? ����>�`���lP[8����P�8`bjW��^��K���I�]q�N����������X �]�T�C�-���R����W(�1�ߦ�!�5��0p/{�_�������Ѵ��@���Q8D�֡�s���ЭmVUOգe[�!���s�j*l���̌3hd�������b����D��@R��L����s3xl�rs@�*��9w�=<���vT/zh�]Au=�̧�%�S�D�,�2;)�x�u:�d��?R�$1'n{���`�!Tł�kv:�kX�jS݉���d���'G����դX�|�|�쵱�����?.�2�,����	����*��A�w�7������x��������hB��Y�CYV�Ʊ�/y	u��h��(�H�^��wbA�"$�ux�;oEP�mr˕�޿�T�z�ͺ��'��r;������}sbi����;��)�'��ӡg�O'}51aa�z�h����1��i�Jn��?��`��FN΁\rh�qi�#��g�u�g�ޯ�ứF����r�}Y�ő�pҊ<'�/�I�ۜCT(�$�9 V���3q�n>�hΓ]a�ɐ�X�����1�yc����S�H�"�*r���c����7�|���'
h�f��9#�����%����ߙ'm=�'V^=~���ۨ��R/	�Ne���h�B��3O�<���I=qަtb�I=g(�
�ol�+�JM�e��}j����N�b�}m��-EG4�#�?(�=��{ƪ�o,�b�����~yC[Y7gg�/�-5�ߦ#\�u#�����
�(�0F"��u��0�-���W�7/󨈗��ă̲X�Uv
����&���UZ������y�J��^5z�V`��<ȼ\qO"yb�
�'D]%�E��0M�ީ%<��	�0���O^�	A�DF-b%{I�M(%&|��+Y�����(a�ե��� F�;>Ѣ�5��G5o诘oP��C�N��j�6�C�D��U�� �n�3sNs*4�p���E�+c��u]�HRid@J�%�d�Y��Š��}��3��2�QI㍓��~V<ܓ'6�+�$Z�\���s��qX� �k*F�H��@�U�Д�mێ�Y�Q���g�GH�c�jQk�k���r��E~��4��@���7z���Х�{�;`Zd���[5�P��|�Wxؕ�W����Ј�˟7,�b���O��/���\��l���y-�������G�H�*���x*v���R�� SVs1����H�NL��ǯ��k���k"ٗT���_��g&6�{��`����\:
5?��m��Ӹ��5�)�އ���U�b#�t���Jo:�W�J�|��KH�´�֢��g����ѷ�9����i:*r��4�W`��ٔ�S�S�zcG������E�����W�7��X!�7�9l��L����ب���FEJ
)��&쓺��q��o�������9S���]|#�C�=[~ř�3�OV���jt��v1�k�m��P�͎�7\b�����uD�����i�6Ð��1e�P!��L�c��y���~��b)�G�͐~5�2Q�q%9���3;/���Y����|"_��5�I�rН X�����.��-efo���8���}DM^K���<:H�:L��ɓ�y�#�Ԕ�IhO����RGv~_�/^����8�7��Rt��d	����J�"iM�B@�O}Z��'�����i��D#.b~�h8^��R.t>Hט�LT�#R��v��A���L#SpO<��Ȉ�#,��1��S�v�l�@Ϻ�6݉-v���w�E2nē�W�ʘI*ur�;������xd}�ct2��q:�j��2�27�C|���T��!N큓M���>�C����A�=\C�L�0T����I �����0���4[G��9�G-� �]�f���|�^FM�������Z�~��^��u���h0��C��se!`�u�F��E$�*�D�طXc�~�����`�C�"k��SR��j)5I$�.�>t�����Ga�K�/t���v�[r[Z��W�l�:uX�u�Ed�R8�IG��B���2�O���yx\j��.N_����q1辗|{��
�����}3L�戟.�~$�P0 �\{sDVa2�2��ѕ�����Y2'�|r�q�+H́�h8���d�m�� Z�~P0$'��{"��8JJ�z��9oʂ��dHJ{����a�ߓ�ؗ#rp!�m����?U��2l�c��c+x\h��v�ɭ��(CQ�y>v%��
_z�ȴ����p��i�6���_ ,[o�Ϙ=��5;���$
h���b�'!��ζ|b�L��aSb�I�3�&�&	8x��v��k3�~e	Ћ�s&N��/_+K�r0Ug`f�^sU�9����O�?K����W�7mZ�{���/�f��}i��?�Iu��p�(>G��y�Ĺp��܆aL�Q��q���o�h�Gsə�<���� ���e6��I���q�JeY·dл�T��H�.�r4��jSB)�k�����CcN�H!�"M%�b��`.�1��CT�ci����-��!"ey~�]�{tQN�E��QRS��6���1d�h0-N^�>��9K@;��q��z#�XT��NPxZ�"��h^�u�J����νU1����9#���f�"h��Rb2�����_����˻++�t��$f����9<���rL��ub�Ռe}ϖ��p8�Q���01&7a� ����"Ǖ����$�Q^�I&���L��	½*�m�e�����}w��4�,���\�D�fPD�|Tu�Q��?��wS�6��z��&Sg�����*����s
���('�c��C��3�6��}d�S�p�XfS~�N�>+����Q L�`��t�y<Ԥ�B���xrd�y	J�l��xb^P��,�RYk^6GEM��[�di1v�5�h�lv�����	5�P��ݩ{��S�e��vU8M�Xi2�.�\V�
ai�w�p����]���b��_���h%�ĹP�7��e}Nݜ՟�^����N���uς>$>w���� �pw,��m��!Z&n%�@�DOD�6qh�":d|��{c�'Μ.paS}Ο�uI�����&�|Ȇ$h9'"�3��h7^U%[��"���_��	N�=���������*���B��˅��Gs�����LL�R�%�J�o�C��Đ�/l�ٚ���p�a7�,D��8�T�/��pg�ݑ�N���	��4��~����R(�f�}����r3-�;U�<��2�ϛ��a�P$�����|� �7%ʽ�H��+5盧�FsJ�!'��u\.=k0�F�l5,͟~������r+�!���u����_9�ZH�>,�</��5#nsJ8��}G����lE3���"(�w�+0�����<<63VM��:ԛK��0��+~V��t��p���R�#I�Y�?�fR�a~=�=�e���)�?�ѥ��:�"��|���G��T�-2S��u����d�z��H��U�� Ff���ȝK��r���@G���� )2�E��v�h������D\jֹFX��1!�����
?Y����$�Xx�/�7���"iX���׎�S}4��S�:��ݎ�4eoM�ϯe'���:�@e�x>H�<IaԨͿ6��;p۫4n�W<i�l�_� {Z�D1z#����K����Jd?�\w��N�u%�$�w<�y�����zj@�j��w$��\C��y�5�]��ê���h'�IT<%-h��v���=l�@W�ܫ�?�J�Z���L_8��F��l2�v䐜�k����V{�|��1����-��s�q�&s�I4E��	�1AP�p���J�򥑸���u��s�vz���p���@OKD? ˛�t6V&�nd%[�_��k ��$%�R�l�Ъ�mi��s��{�s0��*�%sa��A�}�ljU��N5ig���&�r��8S��� V��Pi������e�O{���wwF��L�G��c���#�X{��ʟx�!��fc#�
�]xY�D�/` ��W�g�j�p5�����ӈ@����,�����6��]�|-ٕ(O�sN�޼��[YLl\��G�\%&8��1.v\�GA	�)d�dHQ�D�T��G^��K�1�`ꯏe�i~�,<��:T��f$���,��m5�e��3t�EIR��O�����a
��8x)q8E� J���#4��m*c~�S�C�I8B�ϱ�z���F V��2f��u��
�@�&��V?,f;��F�V�<Q2��5��XV|�˱�~E�zql�= ��	��@�G��rg�j��X�B�<N���y��L:����nU���n5�:U���4�4��WSHݶwa&]G�H\e
}�9A-��2D0�U�ǀc.�@5�2��ﵭG�D=bTJ�6�ȥ��VR�7s�-�-��ķ��:똬��1-�蕞�z;V��FD|��w!)��*��P�%X+���\�J%��	͚���,��$~JK3RݩyC�]Vd�������tFށ�-��w�T����xE���i��K��ݐaV�H ѵ��̜n}GG^M�`,�H
(���g{��F[�V����z��ڬ����ȆlhV@.���u>]U�� �ݡ�υ�����%X��3ѱ�.��֌A���8�FεR�抦F���7�/GRq��E�69`�$�6/�i�����<��q�0������b�E^��<G���W����d���pF�b���z���b�s-ɐ���9��*>�T�/nY`@L���T`L�%��:N?)^��t�����!ԥ�$o����Μ`����F4la
Ȩ�V��5����'��|�W��tBP�C{ڎ�A=�Jy�2(7Wq�ԣ�~�x���a��ճ�b����\N*c�������qP�Ů����w�� ��Q'��`�w(b�^�N���r#U��PYI?���/^�W�\"���C�S,�\:��7M�W�6�8�A�mj�^!���ګ�=��[*��^�D6�qr%O�(��8���%�3|F,���0�Ry]%c[���5X����x���wt���d畮��"�����_�5�@��A������#3�u�R�����8x<�P�*���ڋ�����6j+�b�p�O��V�0���2������W&e���&���8M��F����^�o��Ù�1Ͷ�z�g>A�F�x�����o�飺�A�[�P��ҬC�ܣ��s���۬�0Q�:3���1��W���^��7�uZ�����>{��!��>,4�k��>�Êy���������=��4>!�1k���$��f��,�ev_8�F��8����ٝD�n�i�G_�mHn7b5�)I?����K�I�,�1�F��$��-~R���{��]������{�ǥUǢ$�r��U�O�� �<%w��-_B/�lү���e�X�ANz���'��o3���mF��q�2�U}4��g�9=7�gdfy�1t�ۓC5��V(�?U�n�8�/@R�ࠜ��n�ֱ�v3�~��R<0�;bo���/����ޅ����@��Iؼ<�7���bkN6W�!	\V^���,�2?������-Q���'mǢH�9�1�p�g[�3-Ab���ӷ'������n�7O��s�|Q sꔚ ��������� &F3nt;E@��*������P����|o��+/���J�%<*���s�<���2t���$�i���\�b�9}�;�E���QU��`q��q�1!����FW� ����זw�,ÁJp�e��<�,#�VP�iV8�<�(�h(EQ���Zbذ߄�O-��d	m�?�496&P�~Pw�μ��@���O�i�I*usn��;߅GDO���� 3���	�(,/�T0Ҁօf�~��{XW�Ud��/�v9<�@���dx���p�G,m|+�M�ȏ
���"7���q#˃�����+� lW��%��Ulو�[u�Y:E�Jݵ�h��1�VV1��1��#�M<C]� 5�Q2#��.R�_g�"��9�+�jA�-���#*L|�~N��h�U
�Z�N!�<�_K�+�y��Q;����1|ʟ��V����-�R	�� XU��0�[��GAQ�h�X�����T̋�Ɓi��������5ߨB�� ��������Sq��k�FҜ�EAu�'O�:Z�bo������H���օ�E�8`<F:G�x^�������{:eY��
# &>��g�?;�ě{���E�n+����P���6�
�= ėn�Yy�����E�v]��`�0m�	��/�{D�|�'��ogY�O|�Lx�q���}���[)4�|8�N���y�Zҥ;��vt��{̕�I�,iA8ڢ�6}T-�]���,YV��z}�[Q���Mb7wA50H����5˨���DH����<�O��]4O'W�:��xB$8��]1Ա����J�+T��b1,$8���E�Z�#D��a���F�"����BJz0~w��=�����U�~��N�I���Έ�!&���m�d(L���:,qS?�ɀv���C4��=I��e~#�۫��,.zb9�6m�
p���p�r��ib`� �� ��\��aS����O_1	aN8���ȢU���X� ��Lq���6z�?%��b��Cl��S��2�QD3ҩx9��m���\���:�6]�:]���nyE7!#$F��ՙpi�N{WOv��h	���M:�3�`ʬ�(�u1�=�f��1���
	1}--4A��9�1
�·�@�X��a:u�7�Z�+�\����Mo!�0�!'�AK���-�NxT�"|���0�<�,Y��<r�����P��ؤ�-z�˓,P�����-1�^\Xt:��D0L�uչC��z����דݦ����8;��Q���sL� qoJ31�����,J��ZX��@��Gth�9�?��y���S1�j��a��%đ��pǍ�FD`����	��*U�)�|yI}�|��*w �Y�
���+di�O3����;�!��{��Q�����Y���h]��,y��Ԕ:m������C����Φ�Ն=��%`n]�����0�����,�ָ�=���s|\6L�[�D��^d;�uc���2�: ��9uS�O��|�1/����R�p�Vt7F����+\��Z`�Hl�ݣ�p�qJ�ܽ}�4g��^35��� ��>ԥ���d��.l8��1��eZ����`��V�>p�?��v���Xah�71,�%�����p���Mh��7�e���+Y[�@���j�����8��Xs��(�b�A����rs�Ǧ�^�]��j��E��5�t{dI{�AS6�p���B�/���Y�ZB���g�~����[@�߳�XZ��q�W��0S9��}��TWAkp�U�e��r��B��d.)�*~ơ���/������W˞��(h��>�5�&}�Y��G9�9����F�ԫ_�'m��|}!��:�Թ�bl>ס�r�9�4�w���?��F2q����������9)(��;�]d%T�����ђ7�l�h��\��� 3i�S�����1)x `���H/u6�e��0+ו�u!������hJ~?�V�cE;��W���(5#S�u��*��)����W[�М�ê���t�g��r2'���t�Q�)�Zb�NJِK�m�#A������ͽ`%�V"�DDyJO�|8A	��y�֒�l��eַ�������ʆ�<Jr,~��d�tP��=� <˼���ڜ�T��19Y�>J!<i �Ƹ�Kz�󮆧��j��h����TR�Y��fN)׶�T��
?t
3��_���l�@����k���P#i��b:�����R,I0�ݍA�����fcql�'�}�y��73�Է��L�"�Q2iV�%�!/Y��3[���{�A\ ��ww|*�H)��-���� xkbAb�8T���]sC��ӹ�>% 8�,gMDI>1��sd�$��R �ڐz
����D���3���eW]�4	r��%�k��(�r/9��vI��w,��i�>�>3��SE�JO�D�}�P(9��􌻎v�Wg���61�!�W��c���&����X�J%~��R�Zw%�}1{ �}|�+�%�8�+���7�v�Pr�h[ͅ7���U�;�m�o�J�"�:����N=S/�4LU՗�%2�H�a(�S9�$�n��Q���pu�1���f����f�΃��5���$չa`8�cc!�B�ߛ
��fa�Y���ڢZ߿���#K+z؏���^sb"�*�����"Z'6S�F�^��ǡ�k�8��RƲDO+�Dh�����8�������Wseӏׁ���a�Lv4)���+�w	|�{I�v��$�ҙs��b�})�uA��B�(���=A�z0�r��� m��-u��pI'�u��2�c_E�j-!��ue�W}7�����'7���*�:�A�0[���Fv�<vIz1��>�5K�u;iY�Q�Ǩ�B!.G��R�=�3Jk�WG�H�V|���CKW !H>��;D T����n��R4�����D��D�Ȗ%�,�)<��|)���bZp��Z��=s�<zO��F|)s�t��t�Rn�R;�,�x��Em��oE;�~�"-�i�8c+�WLOb�ߦtV�+dl��a�_UpN�`�8�E�IrBwa�#��0��)�iHn�g�~+n"���oM�/�hXAN���әTFC?�)$;�����5�?��:0 �^��x�@�"�*�0 B��!�#/��ef%��䶶(���j�h���L��w�k��'�)����va޳��~�^Y�PM���cӖn��j4|�O��sM)Si��#ZE�❣k6��'K�ރ�Q�)�8�����h-���/���nPi��w��iaCo���$�u�@���^����@_��qC@L��M?���}h���������T���/���\� �������i()/����09\d�_���݃�2H������r�df��r1	>R��tJ����$5����ǻd8��_Dȋ����Ī����}�U?���	[�n"�t������\�.<l?|�jɡئ_p/'�d"
�t�˭r+b�v�h��r�EC
������2c�d|�v9�
VE�<�V`A.'ʜ��,�(��h���j�˱��
��2��>2*5��NO�����Q��ڨ���+s�����ؘ�ߨ|��mX��!��������O_��%�u	�ܕ�o],�o��7�y��Z���_�Txԓ�P|���K/�1��*��hAu��o�����,n]��aΈ�!��52t��<�.�g�W���G�f�u�۽f�]aƧ��؄<2+��b���ѫi?
5lfN��K9�J�"��Sށ̩���0���9�tDIdDP}�zO�y�5C����"���j\s��:u���7����#e�����k��0�G�]�c#�v�$����L��)��PPLXO���ݪ���q1F(�;�y&�%Q��#�^�R0��:PK�(��������X"�Ϋv�)�I
��A�x��������p�MM1� �H�O`�w��q�q%oW֡�6Lp%)[r-���1�L���x֒��A�}8�|x��Ȏ�^ذ��%���Dg-��QH�32�3DZ	�)M��4Evm��?��+?@�yFQ����.��R�7�O���ܴ��h���o��.Y�� �����Ӻw,��Q:�~+��Q�Q���=d|[�I��	�nJ��6�Fc��;s-��4�h �~¤� wU�۪�c:�T�	`+A�*��{L�q�=�]�P��	 �z�n3��عfs5��>x�?�i�*�N���/dh�n7!�{I4ܺR���I?���[��J�,����T8]m�e��氳�Cװ�×�_帱�����'�8V�z\Y�>oG��fP�x9����S�a�7�t�u����8�V=�A��w�._����jTG'{�;9�;���T����P�c%i$䌕�pQ����Mr��B�O�M8LxK���i���Z�$��X�'����dR,�3���qo��/�{��0X��&��U�An~��V �����ؚf�lf0	 β��b���K�B��f_�Y���y�����w�	���R�F�s��m�ey�ԗra���s���ir3��J��˕=���k�(d�Y$�����Z��>�5�ϥ6--[��H������mL�	p]x *3�mb-�d�.N^�w\]Ý��i������
Nʴ��J"����>;x�$����4m�!S[�g��f��/=a �v�(#�:�����2�7 ^�Me�����/-�v�S4�P}3S�:�nns����5������Ѐ��<n�@��>p=(�ɴ̕l�35�r�1��ą7���@�E���%ңFa�Xx� ��@� ��[��:�1��oq�M����x��Q������vd�3hD�"��K`�V�2�n������f'�t@�d}��&����n'EɆ��Y��h:K 4U�!
(6��iT��HCb�����i�q?U�.4�4w����`��
_e����RR�Q���� ��9��~�'c�^+���:�'�FR%Spy����kM�<�eS��>��
i6�! Q��=�I��b1�_ս�gy��K6A�W�V�U��5�	��(z5�����s�n�n"���ձ��c*%���z��@Y�Ri ���R>)m7��=r�&� p9_E>�}�rղ���$S�*��ٙ���6x6˙T2�G��q���I�69�|\P�#	��:;����7���vͫ#&)zDC<�����)[�E�����P��d�����$�B'��X~�f��~�Hd�Kk%#�P�e�3�ֈa��js��?crk��˫�FUJS��n,M��A�m�l2�#k���%�u�;@׵LB��Y\dY3zع�6�s9�s#@3��'g�?j�vsKȃ���d�6l���yQ��f�(L��|��^������1�{�H����6@.��K�.N3�N�{���+�ɿ�K�T.��SU�Y���WuT ꌘTg�$�a�?���Ƅ��#D��Q+���*����A������.�j��y�oJ6Az���]��FI,P��'0x����S��q�N_O뻰�����5��W�i�FC��R�"�jXp]u��n#��~D����$�"7���a�X�D ���Jߝ�HYS������xI��VkΏg�5�r���n<���R3sҀ�'j9^p��)c^"��B������2"k��8\�Ն�b�+]�;��:%����b��'�Dkd<��G)/�Q�3�����[y�ԁ�`���!Z����K�w�"D	��H��W�����_�jn�R3�6�Tw�<���O^j��Le�w�[���*7��Ck�$�1ſ�_��l o��눚V@E�`�MyqfBp4Ġ�y0^����뀬��K�V�Fv;ٵ.Ȕ	;W�8�H�Cd<��#1����}��+�V��DJ��}~j�b���w�:^_n�o|�)lZ�;��s~�U�ŷ��k2���d�bi�L�q�+�}���^al��7z	C46��e[���S?{DO����l�f��}d��ana;2e~��O���1뫊V�.(��ʾK�A����0�f'��h�O:��{�r���Q¦�/�7N�t���Z�Brm����ǆ��X�
�R�S�?��P���e�y��p����@V�TL�1P�+Y����j{�	�D1b@���?Ĕ����ѝW��o����@��Gf^�D�¿11�w`KJ���6���Nn	��A���Z���Ҳ#{�>Z���x"�j��sO���)�*~K�a*
�À��'�߰?cش��i�f�0 �n9�a�}�ϧ;)�( K��dp㮴����4ͦ�4"h�#���J�u�1{����p��A�yl�Ne!���؉&�4l5�o�8>V�%��!�j�U}���^�����<��,NB ���琳�z$�5�|�����-��tǪ��w��7��㘖N�O�w�x�F��d�<�x.L7戰B7Q��5��+���ʴ�E�Oں��3�"�����>��̵�Igj����*^/�PF��w��W�I�/�n;60{�K���"��t_<Q����^�Ȝ><\��3�q�vK��dO=9ǿ�y't����{�e6�WZ����r>��S��]��hōc��-T�LuؔEa�3�c��_��d'�R��}�`�ӹ"�!�����KlI�M��޸X�?�!��o6I�ݸ`��Ҹ���!,UW��S5�,���r!�����&��Ȧ�wâ�^�B�G�E`���5mm�#��_����fgty����!��5�M�3�	�Z^.|؜�;��"�ɘ�oy��b�0XB��anU8pB�,Q��i�"����$�c�x��=sђљvN;*��w���У��C�VP�W�yd�Oo$.�٨����״T�v�s��࿷�{9[�A`�v���0��l�y_�]#�9��f�:ĉ�N�W��}p �M߿[qOה�C%�F�j���#�̝�c&FV�X5��r"�:$�s����@�!ݐ}�=q�j����bn�(��XN�Y���W�n�흝5q��
~u�YV��d�|0c�*R�VdM�䊘>B�L��řw ��:qAE�ߐ~߫�sʐd����V��ߺ�&�M��94شW<!�P��9lu3u��z�vݫ�m���ƴ�wIq*��lL�0������r3��͡{Q�l:z���:�8�����h���d��{��2:�-���3P�����"�Y�ښ����En�{��S�6�D3̸z��yZ..�E��#Ȉ�t5�x�x�9q�����,y}���D��۹�k������I�vcb�5�X6�6�A�\.�q{M��c���p���KQ@�HM)�5��E��k=��$̪V�֜��qOs�2f��ǈ|��iy��J�I���
�$a��=_����ʕ�ޮ��3�;��M���5?�~EH"��L�w��!e6x#��#S��"���}��6=ֽ�i]i{�[��E�Cf�i� Mp[�ey�#�T�_��F��>�d�H�h�z����#��X���z[ڤ̩�ߘ�����8}��ݭ��Ka���-���gq/�of�	�B��/�BPV�Z"���#?�Ͱ��Жt�T�8c�s*�z�b+��,Я���b�3�c���Nkمy8���XC8�'�͟p�#���/*��j�Q���� ��_нZ+��vZ_R�JZo�7ڶ�����a9�`��B����n�F�_��z����xQ9:@�5MO�_2iBpX�OKk��8>��A�:��yt���C�|=K�di?p�����3)M�e�!>"r<�V�ݑx���l9�]��'�Α�C�@�ət0�c>)PT�8Hc�d����;1� k&�C����J47���hr!cl����ݠ ��sd]���>=bw�쉓	����8쾊Mf�G���K'v&������r�xCB��2�1L|R�L�&~��y��x+m�Y�󑾆[��-ڮή��8S�mU�������d����@n-��Z oe;RB�,4�LtR�=j�.}�+g<�e�_Q��O�1�}":���V��#y���$�|n���j�2J�Sv�ׄv���[�IJ8	t'�N����ݽ�{�j�Wb�Z�t����	�dP**A1h�\F�&U��������>��U �~pxě˷�R+�U� _ �:5�n��P�
edSobݎ��aB':e$��	8��/T��C3���J�4=�*�Nh�tL~���L�1Rթ!��NSK��l�綄_H{B�k��J�cSpT̏��P��;	G
	����:K�5���pr�;ǃƦ�gWd���X�w��!i��H���iZ(4z%�d7�B�����IE?�J���g��S���(��1���I�5QB���f�]�8^��h���TuH~���~��7��
�,B��]����F\B��Ӹk�#1��-����M��A~PR3��I��d�^������,�A�Ց���_sI�#�-�>�'�f�nFj�k�I�3���)q6�����s���
#��-R܎��=��ä�u��f+��).�����{�b��θ���Z�U�琴��<���uD��b��٬�>��w�ۊ=w�>�����-�N"֡�x�[7�����#G/n���8�i%H�{�:�;̪[7��#H]b��Z�fa*�px�����EL��1��5��X*�KK��:������0�J�鋠� 3�@���;֊�7�&�x?D�^r��H���'�*4Y0�u�C�"&�m�>U:�ծJ������*x�#xb�-�p�0���±���W�Pl�<	C��z{�!�/zS����$a�vG�M��-	��g����l����e��W/.7pӧ��
~%� Ξb�wgL���9#��XZW�Ά]>�; <ƹ(�'*�~�W���	u�yͤנ�۳mE�yȉ���ʌ]d3��)��L4���O�>WgAM��5�`�ا<f��� )M�� L+N$ͧ�0�&���!T_�4�C�� ѝ]qJ��D���S�L�����,�|��-�lY+_f�t^�cؐ���:�J��|p^v�\Gю�Q%sº���0�����q�iA0�ݵ(Y�G�zE/l�}�C�W=�0�B�+���B��Z@�`�H��v�P?��R8ɚ�^ҋ8�F�۲���;��?��Y���qύq2xB[�Z�|��~��Zx����/�W��uʔ�5��G)$m�/N3��}�(�t�+����z&啺�G(f�f'�`ݷ_�-;;�«�/Ç�����<�K�<yƤ� Ȃ��xs�X���I�,��n̓`I������(ic����`����%o?§�-�b<�����Pm�"�����^�әD[to�.ǔ�jڒ!��(S5b�pߧ��+���>/t���7��H����^�Z�\�7�H��~9�$�(4[C�|IQYr�v�A���l�ɗ�5�/��W*���(?v���6�"�>C�r4�����tp��psT�Ƽ~���O��E����SW�?�jAxUt2���1��V'��=v���w/� VT
3R���Z���_!#�(n�糆S��Smܾn���P?}��JA+F�8)��S1�p���-1�}p�A�َ��SB���g[)CQ�@��W��;`oQg���H�Ko['�� &bP[r�g4���m��|�����x�-��P�h�6M�sXr�U�(F���V8���|��S�ʊ��Q{-n>��؇x����l+��F6��!���#��_��_}�r��l4�5T`B����R���(rj^����?����Dho7�o��)�����7��aN��&$�@9���������3*8���農7��3�m�e��y�>�%T�>Sy�M�4K!���O�k��va��\�,]w��T%B����o�;>�Z������=�m�7��Lh=+�a֍�I� ~j���V�������L��`"-�w�ܹ�l3y����e����U����b�R�g���l')�Rȿl��v+���\Fb�!��^kI��Sq)���x�?��0�u���/��u|�f�W�T7jr����eՔ����6~��P�=�89<�C{@+�f�,����쀬�0�Z��s�ӗ���It��Ӯ\ƕ׾�cy�1�`�\1I�c�԰�����Tc5-��O��*I����-õe.Fs(����o�5 �G��bV���#����ȩ�u��`���rHQzf�>��'������9�����Vz��ݗ�v>,���%������>u��^�#4�(	`l����H�;�#Нs���$�Ҳ�Qh�L\����+�[�A=��Z�~v#�^��q}G���ud(�ځ$����,צ�Gw�E�\ 0�7t�I>#��`Q���h�xI��/�ɖ�z��"��]��l�X�մ��G��v��6S��觮��9�j�pt�s-Zy�ɪ|I���dO�y6 �/���7ʮ���b��/IV~��vG�� �;ݳ4��i�r���Q`���k�$lBR�r�������ly��Y7���yP��3�N7ޓA���K�b���,�og����Ŏ��K}� >7����'R�oE�S�`qb�m�ڰ�tϭ�`��υ�l�dG>��T��̅ٓF��Oy�[;��R�U�h�L3ñ��/�GY��F��ʗs����2�1�+�߉Y�`i�Ց�Ml] C��.��NCw�dǃ�v2N	f�8���˪N"t���8�DhR����z Uߤk=��3J�����!jMs��&&S�,���<(��h<��pp�a����߉�����S�!t匫���h�׬�����av�� �y��)�cBd�XHE��?MVrB�����
C�	�����'���v�����3�Ж��5*$dq�c�fHE7r7��#4,@��:m}�W�~�]�ԏA���՚d���Oǆ�����i(S���bJ1�&�E���A0��{�O�ف�����yP�@I˃��_�
LP��Fr�
�r/Kz���B���˚͊(�b�w���ue5��V�.P�T���+n9!y=N.�_L�����^qT��<��x�qm(g�Ա$_�oc���S�|�2+p�~���'�����8i���Q�ՙ���Slp����gط�˛�)�[lnO�
9Δe�Z$a�n$ӆ����X6�^-�#]ҧ��������4�w��g
D!��ـ'�x{:ClI��m�pL�QX~��6Y�M���&��=�p�� �UIn�@��R}����@Fcn7i�_	5;�{�3=�/y8l��{GX�*�Ռ����{��y��K��l�ۊp��Y��'���a.�Yuӟ�B0� ϲ�'�ȵ/PCt�*�ڇoc-^�J���Z��տ�܆����i���XL$_B^�$���':?I�d{��d���q�J��ƣt�` �Z�zfv�d�n�(s+O�1���uռl�,3&�X��f$���w�,�©;
��rs �:z�m���ZA��M�w�Hc�D���{��ݎ����`b x���^�&g������I�օ����h�ߵ<��_X�x��_�>�n(F�X�����n�K\%��o��<�h����]sE�K���`�Y��
���K7>z��z�=��B�'�n���+jߠl/R��_Ѣ�jg �D@���x�z��+4İ��r����B��,j�U?���8Tŝ4Is&`+�W�O�LVti֪?'À�l��oY�1G�?�r�?��Gu��I�z|u#���U:9phn�dƲi�ZϜ���{8]x����w||��q��p�ߒ���	�D>�Q�3�ߜ0E4����s���b����K-v����0��ӌ�������]e�)2�2֔���R�K��	�T���̀����"{M t��z�Fp�?�����3]���&���՘����1�}h�����;��n�N����j�I�v�F�t�*'{Z��Z�F2Ez�ע��v�A�[��7�Kim�hn�N���t0��z3���zz��ü�j+l���&��&ئ2"�"Ί�q��.�s(�NJ��͎�[�� >�J ��` ��6���AĤ�v.��{�u}�|Y�F�|~�_)#g�R 6�F�w�-�h�X�����&�;�5
Չ��ocuv��2��v�xr���,�l\NoE��E������t��_Ǧs/a8v�k#r��9߂�y���1�>�2�
[?����9���Ć�� (͘�f�K��L�n�} 咽 ��)�x��}c)ܫ�E��1I
Q���|�F�	�HA�Ee��Bh�y{�~<���OH�-��<h��n�9�60F�.���Q��I�Xk�w��������҉�W>����h�)���^ŀ����j_U�zw��&�;�gG��9����Sw@�����~ڈF��
�p	�Y�Z�b^,�����J��c��kO��6п��Z6���Vв_dF�ڿ|��هk�F.'����ߓj��� �#�Ԅ�f��ð4�P�AQ�5GMj�t���-k�%��I,�V�AM��U��<��5��V��������ɓ{�O�nQ����d��]��D��.��p�8��˧Z:��~���?�'�����-�V�b�T�IU���^���2F�OmH�S>qMݯ.�~5T���X=�秱vn�R�{=9R;�^C=�H{}?�d�ԣ��_�2����Q�+'���C�F�̅vA�E=Z��s�x2�۪!� D�02{þ4��HuߘӒ��j�>�$j��4A���Q�S�Np���N��ꠁ	ʅ�6+n�޳�1�n8J<4��b��� �Y`[SM��dNK�z����Nv�FD��=�U�`e9��cxg_����\ ��tyI��_{����v?<ʮk�Hp��&N5�����4�uZd��o����8^;#�:Zy��g~�,3�t���#����-�A���V	m�}������^Һ�ᆧRip-P��_�a2?�IҸ]�ʏnSR����:(l�<f;oR)z?��Q�&�:���՞��P%�Q�Q�QT6o3��WD����җ]��Dn�unޠ��B]��{����Y�֍pp��,-ר{��X�yng���q8m>~sz�����5�N��hU!oE�b�����!�u���(y����ҵ|�7����%���w�5�<�m�6�^�)�:��] 2r��M-� 
"d�@����W��k����gG'��̜�Z����$g��ef�H�i��a�S@T�Z�J�r1s��~˃)Q�pE�;	��B�~��6a��5a`��׈��f�_z�v ���u���4r)�vs�t����ԣ�y�+�/'4_������ҜU�5`�O�uǔ�O&:�!����&���qӊ{�t�D��=�bo�#R�0�!ֽm���@x����o��%r��s�85L'���"q�X��_����g:�`U���!�%��l�r�VnC���B5�K��� �4a�l7���FC�����+8$������g�"	ypl�����	��y��N�K4mH�y#��E�2��J��K+�Er��1}��o���3)�KP�o̝��b%Z�oE�6�V�j�"^b�<=*3Z:��ͳ���kڨ�SP��3��zig��z�)0��)�.
zB�8á�RN��>we��u?��"s�8�^�H��t!�� V�f�]�����$4Gs��T�Fc;���0�M6���u�$�s�k+��}���m��8�)��.��g�������<{QX�����΁�8�x�Hxu���ޠ���l6G��v'�KR��|�~^z"�k΍Q��uHb���n4�׏}�3n�{G'Q��%�/�\nwD��*�Ɂ_T0�xb�z���=��k.�mU�����O�>��&i]b �߳��z����kV=�.�����ghUG�;�0��o6� ��.�\�57���'+Ƣ���zn������d,q�!/�U����f{�/�D1�$�6���_^��c�W��l�v�佊���H��.���� {h}d^�qҫ��ů���T�Y�KO�I�2����c�G�a���!�xu]��Dy�  ���rBh����D�l̕XI��U��1�B*�+����?;�OC(��[�Y�1����O�.�p4Ī_��
�Y̅�pJ����U��Flz�����?��'	r�������I[���Ұ�6��(�C�8X$���a�p���]z�P��A�%���������M�fU�z���2���m���`�"?�;x9,�(<2-7�F�q��-^�u��H�!�t�O�9(1z$�㓪*$�<t�	�(<]���Z�f�vԒ�:U���5<X���x30��m�u(T�Z����-�<�0���/�W�&��2���E�X�ZA�S��]�F��b~��u���,K���tjT�4�N��I����Gy��5��*;�E��NQ~�7s]��Mf=T�#0�x����r8ގ'x^��V��ڈ�I��B��l��$7C�1gTҝo��ӣ�[������``�f{�T!��f�z	�I5����ކ>m�+��O���	��ų������C�b�9���҄Ux�l�n@����cn߸)|��6HL`'�. ���k����u�������,Vر�(��o�]GJ3 (�m
˂�I����N��pr"���s����b�G�K����	����:*���{�"��j�2˂r=g�]�t["}I~�6�Ƭ��0��,��ƛ��	��k�N���?s���>������A�7p�ѕ�N�e���"c�z`�:���-⼪�H�Z�V��k�B�,s�a�[�*ʥgSE���[l����B���;�l'=�E���cT�g��m����r.5���J��{YI\��r�������-X�j8��zRPa*M7�c�W2����]@bF�<GV�n�R�B�����u���}�o��XԼ���	�z�U!���8w�Fq�A���U(�� #�(�g3p.�#d�����rY��|�	��a�X����4Q�ˉ�C�g�� ����͒�nv��J�ʞ`X��dj��ԵX0���^3Gb�sa�?k7�D$	�8V�,8�Y��.��8�5��_�,����(��
9���͸�����Nr�N�����
�+u�|i����)!�c��,W�ˏf����	t�������X[������K���Y ��hp�I�P�X�L";��;�n�q��шk����y�4���:�bA�W[`K�(Ar�f����Q��*��	:j֎¸|�7��Ɔ֎�ܝ�C���DM$I����7�l�R�%i�\���a�FJ�G�l��cΒ��{5Z21� #2���@?���LD訟%M�����x�6/7�O��B����T�����^WO�\4*� tu�(�|�n��hq�����s���{���n�P�a
�����B�A��K|�/����r�\7��!���M�*���-�d���ycV�> �
ij4�G�F0�֨�W�u�%;eJ��s���qd	z��I��@�2%:d*<��؏�ű�K�HI�g�0K�q��<KV������X�w0��M�wX�#�`���Xb����n$P��ƅ������G����b�Fb�'M5J��z���jk�"�&��#LtYj�Z��v���45�=�l?��|y����*qO���ک�ؤE��ݸ��$��Tk�-���u��U�"�xqt-� �d��p�a�����_+>6{K�uT5�˚�5Z�^��P���)�T�]d=YH���:\/��َ�s�-�����#|����g��!{�21J�D��$!�;^{��-
H�bgJK�N�!z�!K�\�z4��DH ���-��ه8/W���I����X�p ���Ab����7���M��m�I�g�s���V8
�U����˥Er:C����mK������<��*b��ץl�����7�*��K��e�K8�`�)��_Aޤq����*6��
��/~�ۈ ކzFZ!ɏ)��4jFQ�O}��M��	�J��+uS�>鱪yL5,%���Z������$u?�C��id�$Bz��T�uSR�]S|�i�؊'U&�Um!��)�4Z�-�	�#*��V�)���D8�����2�RF��y\��
��h�B$���&H��w&��]������\Ξޞ'�,4S�A�E'bm��1�搅Y�so����:~ܾe���o��y�e&h�������KlhJ��`xۿ0��Kg�����h�A�Cμ��n�Egyroh$��k;�w�tZ�k'��thA�b�?:��^P��*7�8S�{㟓jv�m���BǷ]'YW�lZ`s7���^L���[��@Ӱ͈i�)L�=R�{ʏ����T~��@����G,
�7.w�	�*��vc�4���'�U�s��4�߲J`-��IM�\������@��R��6��y����"D���8z�=M9;���ۿ�ٿ�I�W2����Ơ��yl�86�{.vU`;a�;��*�͓HQ�"��a�0uUJ��~l$��)tbS��,q
*q��̕"��V	�2�I�
0�O���c��h5�� �{`d�r|
�u�ж�1@7��6$(P���E�r�5j��-w���|{�hXo�O|�l��?E ��Ҭ�g������*��&�"9��^@�C̘�lq_I&'����<3�|Gk79z�W�7�2��
����z`kM���2�#FJ8�����&��g*c�:�C[�An��FH��K���n�����y�}�N�����c�%���U��H�-+|��Y����#j�l3�׳�d*�#sc�������.^�Hwc�/?B�S;��z�E�,S()���!z�G�=����[��Ǟs- ��䇭5�r��������P�z2d� ��-U�L�&י�1�s��R�/��u^�a=�g�fX� ��W)��C�! �4�8���C2>!��*=�H@QA(N�i��Q-��k'FBj�Ѝ]��j0|*
�V�,5M98ci�,a��p�Mҋ�Yb�q���Fq���&f5�_?���鑖ݖ��iZfm�pu"��]�[G�
��N�S��\X��,�qWB�+rG˸9�?.Y[ͤ| K���x��$�U�4�,*�}�8ON}���r��U��C�Qk쮼�|@�{���\���P�hꕗ�ޔ��2��zWJg��2��G��g�<��&ڣ=f�P����<�|�b�z�
5�"L���y�J�U��YO��ǫ=��џ�Nw�!�w\�6�4Ю(LL���TN�c�����G��6mz^����m��k�M�;n�������[�wB��?�n�iN.�c�6�YZ�2q�=,�V� �8��y:�A@'��	���u�5��D��A����O��Nd�ث��֮��ݾݧOA�	"�lOz�1�C�A(/mFzN�|��f⌒�5�ɓah�bҟO�f~uv{��HG1�$�r�PӠb}F�5�����0�xi���E�n�������=Ud�ৡO ���b,�H/[���$��hI��&G�<�i��Yu,o�ǖT�!G���2w�`���L/�ے|�\�R�s�ڟ뭲|�Z�������ؗ��?����)��a�/�$4�5�U>b7�ݗ �#�H�s��q��yS)��#�{/UfI?�å���$���k���w0�]$�X�ˢ{=N.�����XHN;��g�n���/å�;ԙK�y&�եn�4���I��A	��������TD�ˑuc�]].)v�-K��􍗓�ě00x�`P[�K/�ɥ���G��9�^�>}�D�7A�<�m�Q��DvE�O��V��
���;�%m��KĆ��#�Y֘:�$�SAbma<�ё�m)ig=���u@� �톩�3����	��ۻ�=��(J��>�_Fh�4��bo��0g�95�Y�&nyZڴ��(��#��.'�r�,���dt���z�����S��2�Ic�P��/�Ef�a��֤��E>���-�_>��k���^�b�'@֫�Zb�cK%u�4s�3��G�Bj�2�i�^}�WE� �}2A!!��1Q"u�@�NX�(��8Aj���{}��ĳJ�%�7��,	Q�U�ԛ>�(��k�N���kO�n��NH���r�k#^�&�a���~K��v����ԟ����iyb(JiL\��M����أ	X&$��E�1�[�Ԗ��9M�`u�������f4�Wce}f�Z��$M6 g8�TĬ�� ������Zj#��Э�n'��lG,FrE)Kb�RWi����Uue��w���
v*]3�W�h��Z[E@A�U{_J�UD��1�Ru�JHl�P��U��mg�0��P��Y��uqo&���Z��a3[��<�x�jsq#Ǘ��U�l$Y�����z�q�G�oh��P$��*'g�dm!#p���/Ȩh�<@��kw/i겣I��3�\)�1}�t�qo�ˠ�KLx��1�a���o	�"��̓��F�>l�B��]}�*���^0����8<�:9�~��-�6!�L?�Ѥ��W'vUoɁ�� (�yͨ��1�Ǝ"��_~�QT������O�Q�׬�7r٦���dF�"�jZ�UC!̠�C��dC������iw�Y�f�\�.�mL�Ǟ�5Qa\!Fx��?�`�ߘ�C�i�b͹���Mm!w^�7��Tj��)<�����p�[�o���0�K�ߚ�B�U�̟X��#�"%n�`&�0��g*�����귿�:%���5�������aE>��t^��m�Db�H&Fwa�n�3�&���==��:����������ŋ�d��{�nu�h��?�^��=�Td�a;8����P�W9���$��)c��c5�,�"�+�q�W�<��6�������^k�Z���u��˖�0OЧPI�S������OC��Y����$UN�A�r|��?w�,8�!�)�	J�
Su�sϹ�_������EY[$=�Q�n����?���'C`��6�&��;b�<� �)$����U�w.��SJӫ\;X']P�O�j��ǵ���|mKg�-y�oM%���yZ�����d?(���8���������(E�	�#(���NU;�ޒ��<�K\��-��g�C6����u���M��;�G!@��5ȧ����'̎O�v�њ��>�>#i���jE1��[�=K5��?�:4(o�=M�x�e�b����1��@ L{ǩx�#r��:oF�O]?�0~E��g&�OD?�Rz���t��E��P��˱.�ni�VP���d K�d�
e�Q�=ws��raY���ޯ����x��"��3֜R��܄����1S�X�
 �h�L������x���h2�'44�
����ϊ��ڔ5Z��vي
����*qC�!I6 b�ʹ�x1X A����|0�}O��!<O�}Tg҉�<�]�-�AKt��2L��߷
��D%+R�	:���U�uO�{;��w�x�DI��N��Һ�F<0ms'��S�/&������<��f��ᓸvb���g$M�1E1dg�p������ Z9h����^�s��M�.(��l�u2�/��	���������#���n���K8D���퐗��Cp�����������l�S�[g0�t pt'D���0iV���ϴr5����@M"�Sr[�����>*@����u4b?�
,ͼ�J��!zyХak�w�*���]�xB�N�袦��(����v��Ȫ�z��d5L����:<dn�m)|��w����� >6�����1�?d�W𐅼���S�Y��U�,�t�l�x���Ie�>l�|K��:�f�Z���C�@�nC�����>���fa#6�nOEM�9��٪���5<�#�{9��3�6V�:靮��V'Rz�J�:���π-�;���/A#�sJ�P2�+�MH��q9kb���˔W��-iSB��q?�#����p���w �%�Y�a��-��7>r��Fc��19m�����l��{a�������v��8�}�D������&=��h�PL!k+����#� DY��Ok-�R="G3�������� 9e��Y��D2�`;����M�؁-�����Pw/�I��zwe_�+ {��V�z�8$�8����I{�Y?:F�Ć�]�l��ۧ�C���؅�
�����\HѠvk�Z��x���Lp�]�']~�vx�@���#�q0:ʢ�t_w2ק�.]�G᪘v��Pt��FFT� ����<=,f��R"D�f�����Q��6�U�/�T*�d�sU�܆ח@�e	�_/�,|�r�vTdk�Č���=�0۲���CM���\��F������^ȶb��&=��^���`���fQ#?��,�s�ⲗ�uaF��w�(����ׅ�jܤ�5�h��.�����;�R�v���������%~b�ߛ��	�E�8Ք�h>��������Z���sָ�w�S����: �p�C�?;F��+L� �U�[R�@��~#ֺ6�����͒ 87(����T\F�f��bE��}T�T���3�yw��{Y,��Ȱ!��zҺ#џ��TB�O-�Ee$N�h]H�g�pˇ��c��WO��E��m�6f�4B�X������^<ķ�x���@?��Ñor���(�r���)x��3�.7�h��gY6�-_��ˏx+�rS��A�ltvZ�0/s��ze��:�@ ��KN߸H�L�).���*,�q�W�t���ֹ����{.~�Zq-�Q�ѽ�,�+(��r��"t����ޏ�`K��[��`����|�߉)�/�N���e�`jkف��M����l�<9<��B�����L2v��G���f�Ȓb�wY~3C���?Y�U� ��l7~�#�:M�]��a���M;cv���V��^�z]R��B�K�*�>����jӾ�h�}���W�]�Hi�TU��y�@��*!1E_~QB��D�N^� �M�w����T(��rx3~���[���5���'E,%�f��	��JS�E���6���\y�Y�z��yhLߋ����y��< ����"�����ⴖB<ԛ>�t*@���%�uR��V��-�C��2�����X�G��`	������[Z���Bȑn�]a��#�}����;@��W�瀨c
�T���&ͳ�Տ,�2�M��U�)����'bu�\%�Ef��C����\�o�����Xş� D.����J����3y��Z�i`���"Jj��{	kX�������a0��݆�������+�Y�#��O09�ak�{k���RR�I�*ڦ8N�h�RL����^�M��B�
R�at��(��t�r�)z4��ke$ĲO�a�C�J�Y뵐}�����uvL�e'\��Z��A���|P<���<�V�u1GU����B�x2������4������36�B ��n�)��lbOƯA(�!Hi���'�����:����°�9�J9�D^ ,�[�)z!��Yk��s��}�Yd8g.���v���� � �s8>�E��rI�Ғ٦[����\[���l�\M����]��bxyc$Ӄ� 	�$q���o�Y�1��@L��|��OPt����kF��5_!u���
B|�ɤ$�%`);ĵ ��e^��E���vΨzA�JF��k�9B�Ρ�]��ߺ �#�f���T�.����ކ�M�7�m�#�Ew��o(��3s&]<0�����^H���)^\�I0����(�fz�T:���Z��F�����s$"�T��;��C�:���ʧB�2��TV���tC�(�̤�ן�f5��1�O}'�t�5D"L��,�6Վ����f��	-��BdsB}|�����%b@�c��W��G�+���H�K֋��� Ѻ����ެ�h��O�ih{�'��d�z^A�v�����w�%�:��I�@�Z;q��5뜰��O�+�y��H��ǛO^sc��[�&��\YcsD7B%���9���<��丌��3eeހlu~_��q�d�Sݴ-��_*��������?Y���1��˼�Zf��JzM 3�8�_�|��������7Taw?�5��Vz(t�8ϒc��`r�~�6�pU�֫���}"��a	����I(�M�3~6���Mų�B��5�Td�M�3x>�q�x2v���1�*�hEL��Rt����#ߒ�L�6H�y����	��_�5�5n�T3��N�d
r�;8v
�l��DZ�Ds ��#Ly��h���x��U%?8�h���yrj=��
��bd۱�9O�j
�=�lZrt0��E�!�$/�"˗��*��S��~^���ރ�qߒ4l>u�Bp��65^}��Osvg򾄏��Ð�>��3=��-�������KM�����bQsȸ�k]E�R"�}�U0|z��Y����y��+
�����A�Wmըy��{�)��W�+�G��=�|(�oR��%cA�~���`�^-�F��AO��a��6�n��)����#?4H9!8	mO��\E�'&�lp�%Fr����T��Z�Ջ���Ae,N	Yb/�(����2T���ُ\���DE[I*�E�c�9S2t	���0���[_�a�n!��耞�����YF^`ܺe�*���_h];��êX�-�;,eDn��"V2AU��[��c�OC�$[d��|�08lOWy��gH�3_�c��3-�>Jh����	R�t*�[O�n��._�ǼS�=� E!�u�*!.�M[dEU}ϗ�Ԃ"�'��ײhX~�v�%����.&|��0�o��f�}�v	M�I,d�|�ZRC�����&מ2>�p�����K�ͧ������q�a
nw�Ǔ�[��ɣ?hF[{N��/NI�6�)6*�$Υ@�d�ŀ�3��P�*��z�+����ݐ��tou���f��p�A{ƌ\���	{�5�����-f�2�?��h�p���\%�.��T��L ,�l^�H &©0�����X�������F#@_ep6O`�LߝR1�i�K|I�K�';W��"�݉4L���h�a��1/	}�c��[6����*G�<z$�Kb�4C�����x!��~c*p���u�Ow;R�ß�*ڤ8���#j���.N��#���X�+xqK�̡��)F*����m���P) =�O�+�v8�h�B��8��׹w�T���X�F�d��B��Wʼ�%n���f�ˡoi�����""���ƻ��O�^sف�ݿ."�|�����/����'U�qdut�kL���tpB�ZG��z8�R���>���ѩE��Ŏ���������'�&�[Y�� �N����ۡ�^z�q��&�ȑ8��|���k=C��;�Q�^��-�eN松U#�N��R��J7�<G��$z~���2f�������zׂ�#�@7�k���@?�OdL�T��˓������sl�@X�XOE�5����<#q��qk9��A�U+ifM�(A��,�k��[yץ����C�%m]�O�R��<��9}��`�9 ��$U�+x�~�Ţ��`2&C��g�������\z��q�?�]-0�h�`��%dd�n�#̶�8�;���i�V�.�՛��ɍ��f�H#��=�..�F
����	x��#޹"�L�Hz��0���)�0֭;п��uZ��/(nokHrϭ�Ⱥat������5�,A�;� �Qw4X�ǂ�W��,� k�pۥ�MF�w�ՌS� W���s�w�?� +���zG�S�Ɖ�C��2�7φ�@���*�9�|���R�e_��t������
n4��^�TT>�4E���`���v�^����οig	'��a�rG
���Ź�@VߥO���f#�*B�7��m��X]͆ �Z���F�!#�o�XEgO��N[E4�֠^/ь{�ӌS¶!�Ѝ!�Et`FD��&�I�=ӝ9����z������h�!*�=5B}mD�c�4�V}�q�in������y��{=�2��ԍ��ɾ�v��Ă�`��m�m2���c���_��̯���"#����~f!O�����]�����i�a����O8hɤN�;�%�����$���g�Wn��� .h�]l,Ub"�%ܝ9]g����=I{���K�y���@ �u�}�Q��k� 8�.B�ј����fȋ��^>1||X��AWsX�q�����c�g�䜼�i�����d�XZ�:&֣��jA��Db)��:���~|��R�,�l�=4�a|���#�=�0��,��v~�=]�T1�_�	�8����D��[Pu���[7��yQ�T��h�4�r�fK�*fR��WT���Pi�Q�\S�O�0���2ts�P8j���	�뎻��6Ŭ��֭���S���ͼ�<E��۫��V��Q�z��e4 x�C8 24ʱ"��ݛl�7l�n��{��y>";�.�#\4�7����&�"v���5�*%� 3.2>��84��g�����e�6`?���~a@�n�3O���R����TV*k4���q���'��;����* Bp[�����E�A��5�B�&a����9{��D���%����|�x}+�܃�ܚ�1c�����F�J�`�S��mF�T0�q���hG�F)N?s���nh+(:�����0ggJ�Ò,lT���_�zW��C����	/��K0E�����hr�9�؍?��0��y��G�"9B�*�~��16�W�� W	aT�:m��(RTN�/�&B�����zb9ώ�)�KmV���~��E\V���@S8�n��'eaF_�W��du�E[-����EDp�|.3��1�k�l�G��M})/���e9�긶�t��:�k����ƣ,`뗰�yo��:lڢx,�Y���>}%��cj����Y��|<s6�АD�9���Ljs���-�xeK?�/��lQ"������59$����t��~kX�ۡ5�T�^�A�����0��6:Q����a>��#F�Ո�v����(1��_g����!ہ����������R1���S��٧|~����m��x���!�Q3[���:g��mn;�ƌ��j^O][����3�S��Y1�>���b*s������NC	2�u�����O^`ܢP0�w�f-a���< a�p`1 	+@!v'&�ڌV���f��kDe������]�fL��(������e��D� ��`�A�s/]��m���{x:f�@����EI��Na�5.2��}�}0�����z��6��c�)��_���uƀӟ�7�P&���Mwxa\�j� ��~���i�0���V����#�dȐ�	ڵu�@���s�M#�vd3�V�3ԏ���o�F�͒�)-�P�D�T%��O��%��������,J�*zg[�K|\CFD^?T�h���8nh�tB#��W��\�� �i���`M�?T�:0QDz���
lն�����^�k\��Ĳ�E�"�Y�
c��u����L����ʲ0��-$����Eg%����4G/w���< �|uL-,<�Y�j�W}��"E�؋7����[�����%'
����Gt��OHaa�pr��+�*k�k�!D���\�� �2���''�?7����<
�3+�<�ؑ�t�C�Rti�I�J[{>����v��q##hG�2��ُ�u8ۭ˿��P��Q�F����!��3<ځWq(gߛ�-��R��������_�jx�g��R�w�Ju|A��-m�V�>��O�����휙�jV�?NM�bw�H���:'Ҁ0��r��~���VJ�\��!+��f�Q]�;���i7b��C#����<��޴�Z����N(q"���<7Á�	4��Q���J�)HH���${��q��+��,���Ŷ"9Oi��X3���%�l?s�~�ւ�P���I�
k�/vR���KŢ#�����J@3)qY�꣺WJn�,�J:��K,/�p���?U�h�r�wR�[��ۙv�z�:�mYm��Ɵˍ���v,�_ם8,�4ș�e�ؙ���)�'�UÑ%_�G�琛Jj�I>SkT]*��D�򬞊#�E�>�L�dp+CVP����Þ�}}�L�;D���Hr�'�c&L3��!�������s���U�c����!�<����8������vW���R��������+���Ų�
'�N��{�W�r1
J�Rx6V#Y�����"�Q�ɟ��*���EJ��(���|f� �#���Y)HCg��}9�,BS~�yC��V�H�6(�baC����"�ڬ l������h-[P�V��	A.�뺲p�=(��U�G��W�Æ�Ʋ�=�i�o��sh\p�f� 5i�T�ݶ���P �҂�?È}Q43�����K(�U�Jhaf8��
�0��(�c� Օ�@���]�9��;��<�la�-��n1�W�r��%�=2� �M�Ŷc1Z�(�
��o�tH
�Sog)?���<�ce<f֕�]�}�6���8�eJ��-�UH�P��Wc.�t���	�k��ct�0���k���8�]2��x�s`��`N�;�J��a?��$�"KB�T#e4
(�9�n�H�y�ŷ�U��ǌ��iMv�#~��,N)y,��¢�+��O�)y�����X�ْ��1��;�?w�D��*nS�L��1�p�C�&0�r,Ai:[rcq��i�.�Q��Z��ZIţ[���n]�a�j(C�+�QX�l��D|��������H���HE�I�	�Q�@ ��,�$��A�_:����N���'#~i��d�B�N@����~̚�vw��Z�;E���"g���K,�c�I'�>�����eU,�]�蹁8r#��x���Uu�s)j�u��C�}�L����a��&��j�.D�9������F���кID��B�͌��@�b�sgR%�m�j�e���U�_��%���H�
�����͹�Yk��zH�O	����|�Ro)ӈ}c�[�ୱ��t���GJ�giCs��͙��|m�T���铖���q���о�y��|{��m����L�����_�b�Յ��P��:=�H�kf��\5xti�J�~���w��>Z�D(�"laL}��P��/�f�:-@��Z�� !�_��"�O\`9���DkU}�s��j���o@ye��Μ�Nl%,�P��0�V�y=�-��Qx�A��]�3?��ϋ�����;��ቦ�Ʀȱɕ��pY��Tw�
:�
_E�.SBe�~�2��$��A�SG�TW�0�C+ǿ9��W(�0�`R|�Dۣ�+t��:��v�C�C�z+���v�_h�%k�ZOP�8��Yy'��L�/9�i:�����K)���jeK1b�R�#}W��T�N�O��^�YMY��T�$輳�@-�t�k�ĳ�������́�\<H��I�ywK���V�@�?+�T̔�H��*˕ۚ�¨1o[�_��ŏHD$�ǔD��c��C�)4��yI�����zx-���n�����>���4G@2��*��4��7l�0���;c���N�DO*	&!5���|��@i����+2/�Ɩk�-1�R���%J��L�����(]��H��;�@�
*d����ϧ�Sjj=�u��$����^u�)�j�|�n閝
�k�23M�9Y�7m��W�Ȥ��f9bЯ��HL��U���ץ��A'6t?�U�=�*��*��ZRr\��������k����'���+�࠿ԋ�oy(ȝe����?�2����(�X���Hc�a��F�e�X������Ͼ�F·V���i䃻Ӗy(57���JJ�����ARJ���>�j珠���	�ov�X��i�O�~piO�洫�N���ˁă؊���
M�&�KDУ��;E��(�ױ	K�X���x�W	L.QA�d�y�/�DX/_�A	��A-8;�U<P7�42m��q�XQ	��!���dK3W]�O�ZDJ�P>�w��rf��2:�n��3"����G�-��㰷�4�0q'B��K3q0]V���[�O㲐.ܫ�.Y@�.3$hĘ���]�t&��&bD�J������!�ͧ��a�+��B�VoOg��M������G�'�i}=e��<��O)bn��k�#Vg�'I�o��c*˵�r�yt�@E{���J�ʧ�������������.^����~�Q��9���� ���0oLY���s��8n��%�2^K&;���9,t#�LЎV��~������i`���V;�F�������V�d2'��ln��J�9�R]�~��	ǲC��!^�=vKwǎu���H�����GFpҐWP���sd�[�1��/�,6~�/�⊧�%��I�f �a	f�A�dˌ5�Q�C���k����VlzS��$d��M���t��"}�7�ڐOMX�0$��d
�ܻ�$���Z�wD9����J��1�XD��L�Ly7�����0g�m~:hI%��aU�f_�j�	>��a`�a0�"��LJX���̤H6��Q6��٫جˇ:�&h����w?���Y�\�f�� 9�k��"`�ZC���N��!)!Q;�f�7-��{�� ������c5�W��}����|��;����*e���f��}�V��0�]�	�1�1_��=�4qt+@��8�rĜ\f[�/���P�&�k��P�뗻���R_Q$��:�$E��v{������ �s�j3邗��l��1�'�
�}��V���P�e9x���4�1o(.��I�.R&�b��d\/]��#o�a>*�xH�[�H�V�Y����	v����\�hc=�5��1W��鎭��\��xt��e��Z�7�%�p�,C�H�u���|����0F�[���@q��}�"�[;�X+l�-x���y��.@�ew	 U.�䄡(0V6�Gz�s�S|c�<�I����\�5�����C��h'I��5�Y^��˲V�ILr�w��N02�l(j� (Kd�n����՝���Kf�*�1Fm/sHYeW����p�x��5OK�G8xL���)�����bze
�ˈ���:��W�U�?��*�Ƃ�4��a࢖Mx��!����Tء���v��!D5G���|����4ke��w c@�-��k�y��E7�M�U`�7�b2p��6��>Q_�ce�.���{����8,�ʃI��?Ȫ���� �� ��M�a��>#��۩\�"������v���b&�:��0Mł�ɧҜ5�5γ����C���;0�	�yo�r"�GNH@d���;�U�c#�D%6��㳌U;]È@���/�;�v&&����� 	�Eh]�Θz��+�G�_p$��0�t`�L��`8]?������<�F�
����F{�ŶZ���y>���Z�H��3F�XP����X�Ĩ�{�!e�G�3z0��tEIٝGYH���df�w��{����	�vQ�#i�@B���F/���{r3�P�]#�EC��J�Ho.u���%D/�� �Z���(� f�к;�����C�+T[t�X��L�l`�?�&���M��*;9%&�ʃ�_����
�|��іVЉ�b��P*b�Y��4i^_ܙ=�[#����#j��2���j����<�����b���g���OT_��ˉpx������QE��av��=�Ï��,,�Y����WO������on��j&��AZ����:�����B�����A�h
{���0��$�d���q�x�IH@�]�٪���W)�_��?�NB�<	��5���&���V�p	>tqW�7d���+d��p�]�0]�S���sr��i@�q�K�͟�>%��x��K�<�"?Ayp����Ͳr�6�F*��3w]��6��8PB"�rv�*�������������Wɏ�®��&�ψDC��A��ﱌ������H(6�O,��(��${a��n���N>q�"?H8 ��0���e���3��<���k�Ә�7+�	���/x���Z&4G�.��:{lijt$�V�} m��%O�:`N˶
Z�]��b,W��Ј�s1�/�����w��+q�O�C��j����k ��/!��) g�%�\l�$���J�֘H��L���Ö1ù)/sl_�X�yHF�7� kES=9ڬa=��G�gjP	��H[�**�P��5q�����O�A��&]����M�}Ѐߟ�t�ⵉ��OO�ф���Ԓ��pjߌ���3��L��<H���E��1�7��3�*W�w��?5\�pGd���X�`��y�v��?��D%5C0o�$���t�ۙ�h���zDi�PXK	8�Ĥ�,8y���� ��h�}hLf�Ֆu�~����!J�'|��A����l?�[�{�\r ��N�?��*@�iT�L|-sQv��h8M�9��E����6j�5:e$f��b�ܔ���oaMo8~���İb� ����;�5\U�x�K�C]w���6�HOq,ʿu����U�b-�v�,4�QG�#��q���H���&2bOMݖc!��aEDS�cbc�gov����")�C�&��4��-7�Kz�*׬0oRG�1�x�k*�8,��� 6APՙxq겢myi#��x*#_~iș.�?�bw#�x�X�AuXʹ=Ⱥ�$�$ֽ[/��L7� (�~��!&q�U�{lɕ�Tv��%n`��A�C��� �=jN�5�n0�.�1�5`���ֆ�U���@��˦�G�����J�W�L��Kqĝr���
� (,�U�2((��ڔuS���ď�s��~�/�f%|O��D�휦�|dH����tDq�2���ǂ����s�KO
7���5 �66��/�P��݌-�K�d���4�F�8{�����T�:����j�2QC;x���r�!�̅#���§L2��Ք��`�&ؗ0�
���hCFeM�R�i���.�1� ��t�&�]�*���l&±�`6S%p~2�2 m��e���n�c���ߵ�>)�_�r$(���2$����ld���uvy�`����3j���a��\�������S����d5�)��¹DY*+�Ĳpx����&1�@� ��W�G,��8��A|�;���T1�N�6%�T���֙�{�O����!�[=n�D�\Xx����٣&�R��7l+����{�)⣉ss��%����Xjp˖��/<�c@'�y���jd�$s?��R�%��ɾ�d�3��K�]-34�&P�0�v���	��e��L���0�0��r�>��B+���W���c1,* ��p�D��E�W�d_�� ��N=������yoy��:���?�-�F��B�C���n�_�4��)�5���pn��oi�I���_��"�a��~gV\V�&>X3mǙM{��q�f伧�ڲ�|Q�I!�!=�H������?ax-��,*׽Cա9��W��c�*�D�C(�5�V�io��A�o
I����.P޿C����G�� ���(LcA�)����&F�3�Y8x`7^2��۵o2b�KǗT����=ޠ�~x+V��	���Z��{��8� �o�$,�ݴʛ_r��VkD�� �/<��2���rk[֎��W1Ә�Ը��@:��p�6��P��Q�bC3rX�y'V��j�@2�}a��	TiJ�2Fl#P���r�JHk
8���<[�s�S��v06�t�A9�� �������a��Z7&�j���kBe����o�;��t_f@��񠹹�[I�dFM]�TQ��Xl�����6�L����jG�1�H��vLڌ�B���'�ߙr.��nQg*�0�^+�nҴ�"���h���kh�^
�Y�ih5z��cȿ)߱�5>U�D��(h�-r��VVg�E����s�~�$(j�Nc�F|~Ќ$l�;}�/1D�ĿB��b�խu#k�G��8�M{4"��E�&�e��^���?�҉�5�-sl�*<\~��vZ�������$Y�@�Y�b�t�W��ෲ,֔t�6��XZ��3�a�Y�I)��[���Ő/f$�����?-}Sfo^ڠbkӽ Kkljl��d׃���vy?�Hw�gUZ	,�UYB:ż�!Ȏn�k��2�U<糘=:�2R0��\eyNr;s~�wr��:��y�$��)\[<��>s;d�����Md��;�,�����hCO>�Qt(o���<4�R���{�G�``�x��!�g��&
֞C�����q���pO��Goc��M��J?�St&N�%�p]xȨ�u�FR�znzMTm�Ɖ�bs,�֣Z��$�[���
��A5���d��{�@~KL,�_����L>��tz�K�1����:��
�1��$�x$���E���jֳQ<e�:�G9th*'������B��2P�hK;�e���	P�T��aC�bk;P$$x�eF�V6Xj�w�ߚ �t|�u�]���)�8R �5ăJ��(hl����g�g��P�-�����w�$��(����S�dU	k��r��t�$P�t��U�E��}���AP�UO=���ė�E_I�^�/����r��ם�'�𷽓q�I����"s�C����@�Hň#_������AE�f+�IEf����V�欣G�h�`"_��8vM@z�ѩp�1��I�~�d��ĩ��4d��Y�EN;9�C�2��NW�trl ��-�aĀ�H6y -m \,��G
F��˒NHiy���T�ոH���A��I
��I�� �?%���#E��$�m%c�<ŋx����n����j�W���#K�ˎ���~�1k9���D���	�������Mͅ�_,`��,Wٛ`R�e��EQ�,U���]�2���EUY$��v�#�R�� ���-J����9c���丠����`�Bu@���:,	��m3;���}�-��$����f'`[�|�k���Qo�
�`���� �2��e��lVP���|�����r3՛ �8'x�p�IO>�S��q�=
Nˤ9�<N��"�Ϥ�&�Q7��`c������d�T���;��� ���H�U'��q�-!_8�]�R���"���ny�p0��țM���BM���7b����=A`�^&~�F1h	��n_J�q {�Gu�Gm���h���|����܀�����z�����9��e2��B���K3r�+���:Yai����h��
%�L���P�����\�Z⁄a�ҲcdgnvkY)z��	s�^¾d�#��	�l����o�9:Q�L]���G��17������0i�_;�J��t9�����p(Q��%w���ü��l�S�)/	k���Y��)I��mEe.mu���@��c|>c������6��+�e͕���Ρ
� ���T�
p�^I�:�,���R��05r��0f�0#Q���j���L�t�o��sf؝���A�_n�'e��I1��BZ��v��ש�#۾�|�O$�˅>��S�$P�O�P�d�����S��"���F �����>��c���t�k[���Hmh� U��?�&�2i<M��6�&jo��h�<�Yq��8Ćc�L�P~�h���3��٤�\l����ҵ�C���Y>-g�=y�B�U-rY�j"zc��H�?�z����mN��O�/^���>����TmvX.H�_@d�y��U����P
Sˤ�w�� ���Š��+�$�S��#��{�uz���؝ >"�Z�~�xi��)�����X%6��9�t�3<`�f'
���4e��t�MB���DE6�#�5U�H#vy?�s�wAoԀ>����_ ͦNx�4B'}��ʄ�D� B������

[�t;�w�tak�ߗ"k�m�'��?�?U�Ь����v�Z
o�����+�\����mY���W�0�2o�2*��p�;_k}�v�?�6M<�k����g�-ĺ��'3�S�9R�%}���5����b�T�/���#w
�.��i�4��?�x=���a�I�����[�o�Hf�����d+�%����#����Ǵ.#�O�C��A+��c��+ţx=k��+T5^��wv�b'���_�U� ��D�U�c�D�BgL�yݍ-�z"ZON�I���R�)�c�8,). ˃�U�Pt�i5|Ci�1��ju&-�Krw�%x�4�t�9s�ҽ-�UCB���)1�H����u�g�f��O$�����.�b�ۂ$B*������O/��M,K`�<K	�/B4���I��#�������5z�kxڍ��m
��{.:�x�?)6�θR���=�Le���'�֢�D"j]�EnV��e5�e�)���1[ѓ��4}"y��{�T��j��m2�5�)��"F(A�K tשq��o#6��p"�6EA1�N�=�G@�-�9T%��+��/N���
���)(�0#m�Ƭ�ǋ}�q��p6x�%�V�x-=C��lGo	q�mbQ����n���dd��+�੽�]@�&d�Y*`q��[K"�����sĪ|�߆_?XsL3.@y&�)��c���
��`f/�YB	���K���O�	���
Y\g;���6�F�T�[���ٛ��n(s-�#�dO^�F�I	7� 
�� �����^J�mc�{3 ��2Rw��D�H���/���(F9Ц�=��qy�1*&����(|��ˬܛ:*ᵊF6w��aLu/�p(�v���W:/ձ��Pfϧ�!P�Y.`��*�}I�k,��䡲H?/Lf6e�!�97����{U�~C����Љu���?V�-:�	JE	:�]%�[�Fa�ѝ�~M ��wJ��&�f�i1	����ݓ=��w�f32����l�VE�+E��ؔ���G�$b*�';s5@�;TU����}h�)l���3Y��N�����������U�8�JI�GY����Вz��C��>x�K���������j���E�JUFM��)�dt+�m�#&Ɗ�k��?��y�-��҂}���ʩ�ߍ7��#��p�_����t�d�ׄ����k�@�0�����2�k
H�����{0r�#�2�6��[[]�sdb;$���>����&���\�\u
��L$�>ƒ�L[&���i��0OG�ev�,�?���bD��զə�')%��U������gD6&��t88�}��n1�3*���5�2��Ȑ���5o�??�b���.~K������Y��m,��&��<my���/���°�jC�$�-��z}Rx�ڴ �G>bΰ�k�+�G�<�����t`����	T�S����0�KRͱ����3�(���/�^�#Nz�>��w!b��^��{��G%�TLͶ��*��]Q�{fx=�G
�� ���/���5҈/9��w�|���Ae�/���K+wD��n�d�@�o2��D�L;��K'�j�M��s������L%"���oc���!���?B �E��ho��|��M����_�8���_I�����4�}�)lڲ�s`�f�?�6�J��J9oK;`Hꧼ�}>�thk�C��fE���\�R����AH�>�vg.-$L}\�#�w�>��H��������?��E�̆Fc��N9ԄgcAq^\
�ݭ�R�ƶ/���8�ݗ��+|��n���Wܴ_GqC6�*Uyw��\��C��^r@�AɒX�e�z7O�������V0ݸ�I���	=���4�r%��Z^��MUȆ5���j��/�H��D�{3��+�����Ayg�T�J��w��C���)F����L�Bo�h������l'���R���l7je��ؒf�a9�����|(�4Q�`�7���L��74��t�7���^�<��;�቗z�Mo9ܦ�5)�Q����*�*�*Q{����Q"�(�
�%{��k�\?�4Iۼ�'|h��|侼��9��0�Q���������E˻O�	͚9@6B$������d�C~�Z���Y:�On��d��������o�Ml��NK=�XI��q����?H������ �~�}&��)݈r�)<�V���w��zТsq���B�RM�K�NH�T�����55e�%s
���P��iĺ��8�Niw|�m�]ƌ3"�����D`fkˈ~���&r�w+�'L�^ĈB
����_�B	���$�sq�%.�s��<n�g�w�`*��lN�[�3�R[ݫ�a=��z�,���8%�7"�=�#T�����v_*T�1�=|��j�F�~�1w��vm	��l�t~�>�L���&)�Y�M5:� O�|W������J`6��ዬ��X�P�Ug�<��m+uA�&]l_h�tv_�v���g��b]Դ����o�J�Q���{��=��2�'�.�\��4Ѷ]&�0��9����d�|��stxنC�����y5#ńuȔ�#���3$_�%�v�������lZ��Y��u�i���������4�4�� ���%�~=��U�.H�	�%�)��W��8��^T��(�g�W���R���nԂ���"�s��B�Y�e%AF�DӀ3���"=����y�	k����ŒtT�h��)-�8f{7J,�F�q(��-�ȭ�CRr�UW����w$Ex#z�����Uu�+(MI�^c�ίpƼ
��
�#���i��N� ���[(���D�Q�ƚ�Q������9.�BTXFB��wi��)$���������lN���O���}�{S�O��������]@�Knُ�Y��T/V6��#P(�;Fn�)&��܈{�|lS��O�8�\�*��!W��-(���*MC�q�s����)0��x��	Z��%Q��
g�Y�/�4���\m�=�����Ƴ��򥒂�
��u����%)�@v\�w9AK/i� ^��9˘��G7N;���]���dB����ibE���{Fc�w�|�O4� �\V?Qe �~
9,���G��a�7#�f�?����5%���u���H�]����[w_\V�H��L���N��aEX)�8FO#�����o��%�;�^&-�����[��7��X��W3z�o�w��t�}�[���K ��pD�jb���Ǚv�C5�V�6�F�cx��8Fݭ�	>���'�Z��Q��r2Җ�\��}�$I���=RtQg**0	���eF���
�)₵��`�Q�� �+��8�^8� ����}*�R��gQ��>�OV�Y�R����#�[1�No���vK����š��1�o��[w��.T[�a�RD�����)vnF��Òkp�+/�$}%A	IIǟe��g�2��B�i z�t�=�p��^�Rk�U.Z��#��&S��,X��-)��ۼѤ���*<@J96$�:����Vv�K��LMK�Y���)�O#az���r������G̠�2o7�P��=p绛Õ���hak�:M�[�o�x�����)-��b����rT/����k��+AO������oT���풚"����% NqD|���ࡢH�-py���a9��eL���,�Du��R�W�-���/*��_�G7�l5���0�����x�XA���	�vǉ��#�FÆ�r6
4GLP�N��yf��_�1I��5n�x�2 �o�]�����Y@�j�&�T^��mem2lY~�{t�{� _b�����
%�W����Gxg�uf�&� Q<y����v5Fn��4��.��ƞ~��af�r;��
��G%��q�%Pd��Q�9d����{�y]��o6�$eՂ�Y|�KJ8O<o�e�ư��x6Nǅba�l��M���m&����Q)6'��O緪���A��U�d��<`96XP�Au��Na#��@.��@+v�� О��Av9���J/g�� ـ�d���,Sn}�-�X���O����9ѵ(k��"i��.�1%�D��Dn?X��GHt��@d3��/��gj�̤౾d'n���֨#�}P'�� ʜ;�(�J����zI魃r)��ss$��G���:��L.E���K�fR,�p.X�9K��e��K��W�����l���K�]���5��d������F���'$��_QԌ��p��pv;t򎏤��)��-�B]#��5�C$�3X�&�}���Xs�͵ �^G�"��$�&��:G�V�\�{�����Gu6�,�U��:�������L�[����qԡU
�AF�(�E��Ζ	)g�ml[zv�l+d�UV�u���̒���� �SyԵ�37|�@���g�L�׊���ԙW��.u7;u8�Q��YG�1�w���8��l*Y �hҧ�q,d҅=B��)[�biB�(A8��iz>����M��d�k�;��ؼv��+E��/�Y��`�.�yE�S��#�O��[��VL �Ko�XjSq�l)U��?h�fA�M��:��i�$�p��֟#�ѝ�Kq�F9-������x]��H�O�`n]���3�ݣta�n�P(r3-޹i樽�h�	�o~�	��ǅ�VS#i&o��}M���Gl�C��+N}}���U�G��p4���Y�˘(Qx�N�z�C�vg��Ӥ�P �'Ob��w?D���sQ�ճ�rN����S�e��'-�N�:���U�öY�Y]�f�!_P V7��D��q���C��?F0�lo"���g��`�!] {���by��}��d�)�m��d�"�Z��@ُ�Xc,�
Gч�����5o��G���L�^�3�T.Sߤ8�����x2��S�ͦ鬞r�w��r�֌��4w�U�<FKs�Ph���G������8����9�~b��LE9gR�r�����h{��K:w�l���;L�ͳ'�2*�/_��~��U.�:�c\��JR�#�6Fɜ�z��Pi��x})v��|�wD����h(�`ƾ��I��˳��.�����V�;%X�E����Y�����E:;��a"o�V���|�Ȇ��Н�yj�.�ړ^GT�g�7el�V�E��ir��f�KD�N�
4���"����W�]�J��ѓ��9�K3��Ȟޙ����^���l�;��6�;^��n�_ ��x�D�L2��/�$�
<��Z|��.�1�q�P)U}���[.5�Xe�M(�N Y{�A�|��C�10.�o�o��g��<�@�b�a+T��a�F������,jN=;��.����ۺ�sdX�+0\�ahYw��Sŗvߥ�|�6������7��$��*��څȂczg9�Ɵ��W����뫔G;]=ݦN���Dqp+S-�'y��0+ɜg������>��gIk�(4����Hm�^<L�c��t�_*f���e�^|�A��B�̵Jy!��=���W�z�ح;�\$y�ZX�����g�G�c��D@�,�սt��
,x6�j�%A���FL�.����5�縡|��l�Z��:��������Z�xb���8��芪�CR��#���}��S��,���r�@1��H��"�sĉ���;��LGY!j=\E��{Q���(8�j�er���ntљ�؉R`�t��q�:hh|w1���Ү2�F���~hM`1K��JY�Qm�V�b-�,N�xk�uW<C�umc��@��W�3ˡ���^K��Dp|���#�%�0��v�r�V/��ީ�̹V�ZW#��NE&��߭u���m�r�#��i�Ӧ���Ճue�±�E�M.:���)��]��x|�lCT�~�Y�L6�Mc,*�G��Х��_�b~_����e��-w��p�m*�n�>���tR�;��E�e<$����3���y���mӇ�2;#6�I��4'��lΏ�
��YX�}B�:h�h-w㪝�J��'Wf��O/Y���Ez;��( ���3�W��,�֡b�ʲ!���è	�c����y�JR/3e�h,`μ��aKg�d��~�ڂ$K�)�V��F��=;���Ű�A����l ����2[��, �L��]jP	�i����E\n}$F#D�\��:�vw+Z=�f1���ŨYP[����y�ݜOƷp����r9���Q�O4�8����'<w�?�T�N �v# ^h2e�9���$q��y�!���v��� 6z6_jRs��d��w���_��@���w����'��].���!���]O`y%c}������v�f.#�$$�/ց���ݺ�$�O���~=I��/�]������C"���tE�K~O��0ԅG(n��i���Q��-wey� 5���� �K�D|�'�{�x�R�m.�O
�{�(��������Z��6�"Y�v��q	?!��t=���>%��n�R���U�ǭ�E����$�Ni��i}�v����eؾ�BQ}���
��t���p���Ź. ��b�va�'���n�ln3
�u��B㴪�Kd�50R߬_��tOG-m �͂(�J#XV�@�r͏(m�c��żި�^��������d�9�� ��b�0Κ�g�v=R���{��@�6�1��ȳ�Fe�t��t��_YXr]�׶i2?\�����h�_�݆��^����G�8��:4����ϥ �t ��x8���-9������
�h��E�&.��دڂ��9����k�E�r"���n����5���=�� �X$ۅ�k��f�_��L5�Q|r'p9�b�ZE��ӱ�C9�<�u���HN�O���hU���8�����^}x����=�ԡVwt�2E5��.�A��˵���G���:��+2�����k�8�1�.?o8��`�%��+ģ���1�+*ff~ʅ*��[>�@2a��������N��0��!q���D�D�KW# 5�=�K����|]��+^������y4ݵ�=�؛&{ܞw�S-{/�4��l7wiXьp`���ǯ�Bl��+q@��}�����'��iy0��:<�
7ƻ��H]�/��:!�4٬�;`,?DR��-�:շW�/���3����=%b�'�1�-�
VC|qm���+b��s��[=`B�_����U��� �&�c'1Y*��{ <�u���AŇ�t��q���Z��VW��"~��'iD1���+÷	��+����eM�������:;0�ڨe@^<�Z@�)�Э�kV�4�|�߰��y�x�_3K2{*�Pb���Vl����pő��Л��$������a5�ؘ.���L;�!��~�tR�5u��F�1�6��si��`1��9�/DK�p{k���O^(g�nlK��j��B�Zv���F=��Ow�.5>�
A�ڢ�6ͩ���ы�$@pPTn����9p�v���Ӣ��2�������u�x���.'F��ȵ��S3b�1b9�>��3��!5�"�o��8 o�e6��o��opK��O�0{�ʝ���ww/*��&j�H����%{��u�^�,���U��O��ъ����"���W0��՞Br��ۼ ܊aNӫ�$wEß�`���`zc}���-U�x � m놂p���m��M�B}/���)c1�7J9����/]�:5�Tt�)����G���*6z�ٶ��-)��p��o��x��،�Ɩځ���y����[��!(���D��:z�V5�o<i^�:Ї�5�1`��b����r�ǎ��"������;,���x�Zy½l ���ь���5��c	�>�(��e��Y��60eEQ�A��Ҝ��c������O��%����'$�:/�j
��/��V�O�mƇS��?��2��vl4XAIn��t���J�(�(�F�pLT WJX��~�G;�krs}Ƈ�4��p�D�<�(("��q��W*�N��ǀ|���z�Ӱ�~$D�1
��J[�}��^�[֬Y��fi�X����Ik�b«3v�1$������w����A �+-��>¶h��\�;�DRe>����xTJ��ѸFi�L�R�k�Yj�!٠*�Q�W';��{�utoy��Uji�5x���Q����J���tƟn�5%ǌ�7b�z�:9O�Lr� I!�2�D�ۡ�*�@1��93Ah��r{��9 ,��q�x���c����Zt|+�v�>���[�s��3��U���5��` &�����)Iq�=�����K)W��>�=<��̄�ҥ� �03���ex���b1�I��+5.��Ǳq��Yg,�1��*��)�j��! �|������Y�ߧ�eV?u��4�eG��
���9 �p�{Gd��X� �\���(q��=o�?�U�L]�!;��t�ź�?V�^���ˈ:T��O�R[�x��:��L��b>QWϨ]�Lli�PpƟw�W��>�js�Yx

�&�*?��6��/���ӥ�8G�
�06үÉ�#�#6|��ИC���+΍,N�ro�u�V�fW���j�sݳ�����ON��0H�%�i�v�`��{�z��˩uƯ�&���I��Ӹ!��tZ8~j�ji�����VH� ��o�l?�� C�˒�᭯h֔��#�CNSO+���D��Yk��R�Tʾ�>�J�b�Ή{�1j#�l��~�X�![��0���?gnqv����E�<<Bg����D`@1�P����!�Ѣ��3��fo&�B�����熗��䞋3�;J�f���^骊�C�;<4��}�3��z�$���76UG��q4z�� ��uP�B��Nؙ�^�Gs~a�r�Hȍ�r��KQ�A(����1�%���g�Jf5�T�U��, ��������H'�_䬙�:8UV(u��[HD����q�j�FD�d�F��+7�J���=�`7���a�U�2DX[I����tx����2���=�8VM���a�=c5���{O�b%#/�;�pxb����|����_�V\s�䔴�oN�O(��`Dq=4�����]'P)��ӽi�Ye��Q8\='��!O/�T�^�c�)�j�ѓtdRD�X�����}��2g���1�"aU�Lc��}"Xj�Ʌh���z;S��� �����y�H���v�>��&�J�Y�-�ך�K�.O������͏�N(5�;b�n���8��j-�N�MC�R�g��qnh��U���#�߽��0�42�*�\곏0a�lQm���r,�T�֦_-�G"�7�o;���a{�����#2��tq��4�W�"�prH���3��ѝҸ{�| ���v��,J��n��vP{� (��ԬQ����'pJ����s��S��/=H�U�)S��>�5c� ���������ӯ����k��S��r�E2��M}����Z�@�5�Ñ��F熍������v��������Hci�"Z��e�?�l�Mz�ץ�>��L��
���(�E��v��aV��V"pEʣ�`�������FQ��;�q�p�%��&]��޳2��p�8�4>�$��=@.c�D����XC5z���P���)��i�!�F>�ϭ�קƇ�1|�.��`�3I�KѨO���"�~Je;���T5�20��݇�v��s���g'�c�k�������B���ũWζ��X�����n��4m3�~�5��%�C3k�<ז��`��Ex��}��a��|)�JI�)5�:����q�-�X��{{.��9".S�����k����Rkm��ot������Q��J]�um���Ώv^��dc��q�j�E^�zoK
�F���He
���X��R 0���H��*�|{R1r���%=kbO�@+�t�A6M�H�"�Ŕ
wF&k�ӟ��+�I|ދO۬��vTʣ >"�B�����Nc
r	~�0ҙdm�@dئa�S`�^{��-�_Y��n&7�2K�2��g�s+�d7��Gl��&N�MO@K����W�Ң�Y~��L9�7�ּ��3�h�������o����Zn@��K�s|��>��ғ���;�ᯛ��nkC�N��X-N�F��0%���9�֙�FS�%� ��ꇨFit-�h�|�M��Z>��U�=!���y���3$�ѩ�P��[ܖ�͸o&�?/T F��~��H�剄zVOs	 ��q-�.�2�h���5��]iH�q;���̦�&Y	���]�z���x��-!��ߓ���	�"PXQZB���8şb陞�����xLA+��I�X��{�ǚ��c:��Mc�n7���ҏ^9�X񈌋V�$ �R���S���ᠧ���G�>��!��C���3�V�/kδ�Mm�^������y4w��*�����頣�$���	������~d��ڣwb���&(Bܰj���S`�I����G��#t{ga���4,��=��g�B5�Piv��[;UEd؛���&�n��&���u���~�&K�=�:�&q�_��.zӹJg["�<L��or���C	5�{�U 	2�+��,>�pp]t�]�$�w��HV_�����}�.@�[�|�Lm?5��\���G��p`�-��i�,(�a�@���^�Ҧ�1]��$�Job�h����&����G�X�fr�q6,aR��wȽG���y��P.�S��P�_}�:(l��5���+qwq� ��^��?�խ�:l��+������1��p`��VlF�u���Q�ܲ5�=C/��ۄ��º��|<��)���d���\CO��+3o1Hk��i!W1�6V��S�)�<D�1R�\
�Lq�0����U�ř����\�슉�L ������T�15o�A\��1��U\('�S�`�`��(��D1�'�ys�L[Mm3��࣫G����2�nʟZ���M���{�j��4�H:��%�	�*�2��?������2%8@����=���s9w�G��~��#�����l���ٺQ;b������������@�s��pJ����T}=���<m�+	c��R�t�yq�i�m
~10�|7d@�^�ҠP,j�6�sj�_���EZ���uX�ȕ_�����,��z�h	D�\�8�;�[���?�ljSpe�&�����Z�Bv���naL���7�MVI�-v�*�0�l��j�]e��ث ��V���,��.94�ɔ�q��~Ӹd����m�!S6T~���uZ}4&��L���d�XF��9�,���)���Ȣ�= ��H�x6��3�-���w��S;TG� �8��ܭ�����Q�S�MO���<�G��f���׭���:�ڡ8Ϝ�A#�e�y��z�]��r��e�n�VF���+��3"Clj����CU�/��hTW�gMR!��շ}2��rSy.�����Jvq�0��裣q�f���ݨ�@��23��ٰ;�z=�A�hɓא�>3Q�d#��d�'<ơM�~<w?&��XN�G��k:F�a�$�fx01�cيu5.�܍.��C�y��24U�t4�!*3���b�
cՓ�(/Z*)�����W�v�T��R�=%*@���;do��[����%w�{ͪ���9��/Y��b�������C�,�t&����[��NC%	�5�Up1I'������Z]�4�D_��ٿe����Qgl�j�o��7�N�9z� �SMA:��P'�p��g87��b
p����'�E�џ���(���Ia�۝�l����'�#�5���"vb5�QQ��� Za�M�ij�|GOx���-P@q鎩<S��D�q9� :`/��~y����������SH�=�Z��tj����1�`�Gq������;��&����;,��! �SI�l<�֡�Cԗ!�%B�*��h����v����(9�{oǶ�^{%H<�6��$W�m�[�AH\�A�\2H�X��=(X'�b�9

q��:�����2
�"U� <�`�ϙ��|7�ʷS�8��A����FSKL��s*���1f��?m�p>��P� :BQ��6�3_D�l��G�F�1��%dZ�z�!�؏O��l2ެ���b,���Q?�����n�b;�C��r�2PM>��y&a ��͚ؼ�ݲ�y����u�����i��y0BADf���R�C����[�"��R�����Aކ�p���?�D��?-��FO�:Z��t�G��@N���58���d��V�C��c�r!����/\�5�˟mE?���u��$���NS4q�ڎ/n<C�zF( ����B�+lY�0K��c���o����������/�a����GͰ*�x�ie��e�b�{���z�9@b�X2�0U�P��Ì!�>�-�nx+�>?�5��5[���&�+�b�%a������^�����IBԦ~��T<���GX�Qv<Z��&��{jS����k��%�e�KU�u��+ҽ6���6Ss%_�Cd�L�*�JtN����p%cEU�0w�~_,RI���@����$k�ũ��&���#���9��@:(�s^�LN,y�F"Y_�&f�=��W�%U�	rQ�Vr b���ȶ%�"vC�h�q�o_0`�~�U�qW����#���5�'j6���ۑ���M�i���A�RjHq���ue]o��G������.3��ʜ&A�����>Ml:4p�09}�N�սx$��������Ղ)�z���&�̪p��;G�S��y�d��`fHE��©�
OV�#1�ߊ�8���Q�-��=JJo��v��Fd�����'��g@����h> ����U�{��(-��",��{���t�w�}&��4^�����w�[��!,�����3a��4f�u�xA�Ig��B��nc�,*���84�Cv纴~07^}���b^v�g�
��(����#_4M�>���X�I��+G�%��&���l�JQd-Z؇��1����`*�Q��d�f�Á�Y	޻��,�<s�5%m_'��ٲq��P+x;8�E�c�%�X,0��̺��U9��K�!B��0Q�@��-�ڊ�4��T��U[���hܘ�`A ����˵�x�_̪k	��z`8L������\��T�7��_�����:7�0�b����5�g_,�3�E�6}�"bx���^�I�{���bf��
���j˖�p�!�e63�Z�D�t�� �����Q^?48����T'���ڝ��WKu[��ņ�����<��R���b�C'Gի	~z�;���B��J��҄i;f$N�t�乯ٔa�O����S�J�Td}o���J����]�	�&,�Xs�?IVl���(�Z4w�C��	~�f�cf�,����ݞ�w�<�cw���*�3��
W:ТБ���xV�ח�/��D��,��X���4��;b!b�'�7b���<��&tAƘ������p.�zP�.w���C�d�����3�j�~Hm�\4p�YY�_����"P��=Y�gIq�Ds�,�a��6�Y��\>�Q$e�B�� i%� &յe�)3��*aZ�J\��z�@$�@��H~�	��]�꾥�d��C����nKόfh�⟅5��X���ߨ	�X������GMiTV�������O��)�o����Ƚyd>���&�H�z8�$x)��t*e��yZm[�O#� ^�}Ϸ>�1GU,���+YniA\�	t^����t�]�(`oҤŬ+�dW�3*�u)�B��T����ͽ��NX&�S�� 8h5�،��H�J�=$�R�!O!,�`�M9�>�Z?�_p}2�\��u>xi�x�^�s���I�`hRm�Cg}�g��ͩ�b�N�I��h�烎,��+5�
˦k A��CL�1��^����9	�5F�%%��v��8'�=궾Y�"�2+@/FjA>*��@�R;�z)�s���כ��Ņ���zפ�8�P��SK� ��=CG�oSR���w�8}�N#�i�[���RX~3Hr���"!��E��_4K6���*K?D�!$�So���GUUR�X�/��N���o=n�ǎ$r���I^����9
I(��S��;;,K�pH���~����X2��C|-%�c�-�DR��_\"�y(�tw���!�\��UY��F݌�9�#�yf/],t�z���g��G}JF.d�$���E��Jea����όO�Z���~���
��e��Q,\��o��u�~���O'EY�1?�:�Sa�#�|��O:s$�@ .�[�*�MYP�(Ĭ³����$��z⸾a9눂B߭h��y�k����W�7(UEtoܴ��ڎ�*E��K���;�����ސ�q��.?��Rd-z������/�rL��*�������f˓���y>�G/u����#
�+��?v����4o�VқHS���4���P@4|�Q	<`��i(�{X�M_�2@�}�
���+�[+�H�5�����B��%�I���X!�tB�C���qxҬ�j0�O���M�3I���gu�րH�3�C�c8�W� ����x��j����Ю�w��M��:��M�ڽ