��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V��v�8�fOIY�wǇ�U���^8=��r?�g��[t��h�$ئ^Ž1���/,<:���S���N�)� �$����u��ɒuޑ	�.9dTg����n�Rg�ơ�*s#4@�k���$�;�Y��Hi<�������mĉF����ɢN��A(��<����s�}��E砹{;(���s�	�a���E�J6��S����~�|-or�� ���?w���h��S_}GKj5{ ��n�Zi���W�����	?�k�kʫ����;lk���@�	X��{���e��t��G�'���g��~��M$��u.��+��~���95�Њ@� ���P�HP	�"M0�)Gp;&���>�¼�ޓ< ��ݧ���u�J�k$A]��~)m������1܂�6&Rԝ��,+q��̩_W1�<`K�F���q4M�E�i}����	��ђĤ�0t�w��b�;��;��hӴ�tIp��ͼb�,~ν����/hl�a���g�;8:a���`>��օ��ˢ����{x_]S�/��R�`!�^�믮��*���Sn)���a�/,�9ޟO n��"'N���)߈T��gnf��<2�g�����r�Z�F̌]��!�ӕA��.׈ezH)������I'ԙˊ��64�7�V��M�=�_�o���,q�'^>F�g�L�MVW�7x�����Ju���$�t��v7����Ӹ��_��W�c���#�Y��ܰf�GP��y�}�<2��g	 Z�X��/�Y�Q����"	���׊g��ga%%t��cՎ?��}U_Tv��+&DbϜ�c�������.��T�<J6m+�]퇶�
;�>E�?T�3��/��&(����2�Qwe/B�<�rQ��ei�X��0�������tB�cO����wʎ��e�i�9�}{�'q����t��`�ؐ��Ow��`�7� �A����HЦG����Hõ�yQԴbc�q��ʰ�J5�vΗzϯ���,�'�37�Sy�~�{?@��4��S4�Z�ob<80���S�I6�+���^�<�IJ��i>
=	�y��xr1�a;yQk��%^4�^jZ�E�*�aH �#��bH�m1����ܛnS�zv=z���l@B�t8��?N���R���i%��K�G넡M`�S������}T����}�`�ȆX��vf��sU[��� ��R�(*���F-�/���f"s˄'���N�q�Ж�|Q�t�Iɠ�i��W�'�:����'��Ǌ��=Ҧnls��5s�K�Sn}��(to�h�w�z���}5w2V�Ti��{���bv������aJB��=?cwz�V����k&�E�Y*0Ho�U�"�p}��*���k��-ϛ{�a��-�I�F�2�	I����P)4t�R\�z`X�v>�ѷI��0mf�-�`j���>���p��Ww�i��I��"�W����K#�J�w����L�Z�CXƆX$=f����tv:͂`Fw���a�Rp���t�aa���W�<
�,M@�C)1�u�P*��<���j�m@ˈS|�1�T������q��d����dL��t�$[.u-%p�BP��`	�un2m��]B�(2{�c��)l�o��a���}ҎO���BnA�N?Xf��s|暍��P�_��x�]��/ ���v}j|���T�ڬΈ�vga娯h*��w/��"�;=u��}�!V��|ΕJ�t��}O2Zíu�rh�R?v�������l��ձ�,���N�Y���YhAE�#�g�A�IE�y���;���O!`�~]�k��Z�EDj�����y�cva2�}3�B���spZ�$բM�8$����^`�P�ۘ@&��2��ת������N�_F�\�U��G�8��/����@H4V_:N��z�-���\��s\â��\�g�o�k�b�H��[��VN��w�2���A G��<:]��h�9ϬF��wu�XKs�W=E&�RE��|���3 �>�Hŀ1�� kA.#�vt�}6Jv�b�v�FP!���S`J�-��5�;�8�� o1z|G]�3���z�����~i��#�M�f�q��T�K�u���S�����ii�0��=+���2�l�\Tx�~zVz��X�Ե�@C%�I