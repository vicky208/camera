��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:_f������د�1�Ty ^��D|��K-�a=�����[+�͌�(G��Ɇ������?O)^�� ���$X�ğ�wH�
PZw�/�s����x�<>�"f�7�@8O�Ǖ�f�[�T�*�!H@͹Z�$�����NF\p"� $��̈v�@B�!T;�2+w��`����"a~ӕO�)Y�����k�Y��7�`��K(;Pѹ�<��񁅪C�u\�	3=H!O���gc�nr� 㵌��d��T��D�W:��H/� fn�%$�*I)2��L��f��ppf�0x|��>���0v�I��"��o���//�*U�ڪ'(tM~�t,l]��P���%'�	��|&�}��j��:
ݼ6S �5���}t��r���y�����SI^�~-Y����3ׄl �HԂ�n�z�|u�6�8��c�������J�����ӑ��<F��pQ�"��eA��|�8���)�[ ��)�lȲ=6�~��T���።hw�ȍ�,
Pv�JU7��WB�q�����C����b����r�onь'��|�u�`$�V�Kց��.k/����1��*�^:\_"R���{�į��S��ҵ׊�FQ�C���KEP"o�h�im�w�����e�ߤG��	A`�fۄ�-�JM�C8�1���8�tE��秉��]��B?�F�f�g���Pp��m��3��!!8�o�f�����&�+�:��t]RT��a�&���|cߞq��N����T���|��6��� �}݌jL-|��I����z��ԯ�)K�Z����\m2-	�hL��V.<����F�����Q}��I?{�O��1>=�>]�+5N}����N ��E<��V�n������y�Be�c��h׼Ӛ�VV	e�c�U;���
��*$X�����t{����>�6	�ѐ-O%��bt���2f�d��6������)*;sh�l�@�	��U� �;�o�a%��#�e�#B��>�N�鈸�F�&]m�0x��T/P���**3*Gf��>��K�@�OL7�#��s����<�3Hr_�}�uɥ Ĳ��_��:g��[y�h>�-tw�˨�F.�v��1����U�6�O��6LQx�]��9���f��\�^�rqa�B�d����Mw��[WS����٫�4�X�7�u� �n��=  C��'ttя�{�ܠ��
N�Lo(\�}�	 �f�4��>*�3f�mCb��u!���h�������'c)��ry)n�Rx� ���ܜ�4���Eu�=~.V�pV'�k����ϖ����]cS��Ef�m���!���G7%�yCZ:[���M0��E$W��j��1퍟7�����L�8;�gE3�ȡ��u��!�n��%����bu<���0c�&�k�*�1���A0�n�l�Hw��H�x�:3qT�t��AϦX���->&�w�,��pb����U+��'����3��L�4���	B%]p�� :4����p�����+_1�`��6����v^��bV>�D0Z%ȴ��=�_x���G�n(?XW%θ�	�%Ph�gj�x_�1唋�е�e��4���#��pb⋦P;'p��#ﭜGB�بpދ}�d���r�3�Pmk�<T �IQZ#���m����-����L���U���S��ߏs��WB;���qw���m�����C��p��HiI?�4�둟�g� ���~�Z~�N*<ۉ���z��e���>�+��턓�n�5��5��x��8�0�J�6(Ϡ��b��?�+�/�n~t�f����Io�/��+ǛÅ2	E|��� ��=z�V,�惈�Nc���L�S�EBS�v|����ʙXL6����N.�³�z��2���R�>ZMFBn�'��
Ҡ�PQLdern�?�89��8ΫT�0��Лd�F�x.O~��3��Y.J��C7ᘥ�i$�UNC��U��!�����4=������ؠ(p�'"���N�Ջ�����̓�J��en1�عZhT.��;և|kJHQ�%)(��i�� ��i�,���R{�DF��[ALH��6�$��K�m4��fR�s5L7
��+����	j���]/?��>�rr�!��c�"b`�Fp�kh5i�I oC�����$��YG���5�Ā�9U�1�s��u�꽲]�!o)`��ͣ�oͻ�P�A�������q�^�e<�B(˓L��j����Xk��}�VW` ���m���Ȉ@��3�v)5��3g��+H@�)t���J詒��!T��F�=��k"�˛�#��@`�y���r����p`��u$$�������rQXM�Nq��?��ݳ�Z;e���ꄕ�M$g��-���R�&ыN?D=��x��HmV�wLhab�bBqI ��	����ؾ?�$8���p�{M�,e|��@6�R��
+?Ə�����'�=��8.��cL�>M�N������ iaK��T�4����q�>���8�L����ؙr��������&Sc�pJ���_��΁����M���K�_N�Y������*cE����8֞KR���QrOj0Ȝ"�c�5j���j�ѩ1G˰ZM��!>���
���W�r�!`�0������x�5�����1s�d�����L��^ܰ|)9���>ʹ:*�8��j,4eY��ChS�����2<�W-�Y��
�"�75�4���q�Fk�@�b*�����4��/����ǎپ���ST�el5��ѝ�ƶ�7P�p�B )�I�S<a����[���\2]~?���ϔ�V�+�Z�L��Kfިh���岅��Z��-aj\؎�A˕����pس��'�`bA�D'�W�g g� �ڨ�,���
Z�oK,Xr���=7���-7h��HS��]�-4��'ĉֳ7���oZ���>�c�SZ܃1qYēl�jND-=�l����˧�,%���pDU�'檘ƳL���"Yy�ti>%�y�yq����7���*�������r�! 6~�ӊ��G}��ڬ���r.Ӱ|��N�E����A�{��?�P?W����nt��c�_7s�Z#���1�&H��Y���!$y���bؔ�p���,{�k�a["�����{�FEq�\�pt���y�i���I��c�����	�Q�?K3!HO���0�#���B�h6��`�Ch4\ϖ1��J��,j�4YP��]K�8i��g(�DR�Ӆ�m�#ߧ��1���9U:2C<x|�G���ԅɶ�q<�NLk��	��oL��{�O,��d@���Na�#��aӸ���o2�����>���"��f�h����F�(�їŪ�ع��r3�]'�������$9:p9R�[�R��� @f�c��l��Y�o�����}�0n����c�`��{��!0��@�*�WXi�hA�ʦĐ�!�&������I�J*��U��
�X��c@���2X��fɢJ⎒w�.XKv��{�<�A�x�P ~�����Qܯu�Tod�3~��Y���=Fr��f���8��.����~���Q�}�+��l>�]���"�׋�atޏK�`I�Cאx@O����,>ܹ�Ul�
��*~�J(X���,�*.Aͯ�[X��Ї=ѯ	�e��2[����0���m�<Rޝ�⊖�Tv�7���2ɉO�qR%Y�ƳҺ���.tZ�$������]�%\��c�R,����'�OoQ�u���P(�y��_��o��I�{������KM����ay�g��
gWl5k`?$۵ұ6�]������ROD�W���L�rhz�G[Ȗ���9�^h�o�D�75�1E,�����x?X	�1�.�!�m8h��9`b��Q?Cq��g�-�/"�3�7i�L��oƛ����
1������^��\e�3���]ZOS�[����?("F�W�A)8E�<ҿ��r�Y3�&C���S���d,*�F��ڪ�c�1H5�3vvi�L���9���k�1Q���mR��K��ܫq���t���)[?���+�L[��ɀ�&���+�Ы���l�t�2�sֵ�z��KS�9�eW|�bO�O<c�X�|/Ŗ�w��7q�S�%,j�5\kiܒ���iKK��ʊgW;��v;�ַ>�KF��J�*��6m����:C�HP�|����V�*����^�@ajp!q�C�w�Z�ob���9!FYv��P��vU|34�S�����o�T�|�剜��j4�xנj�����o�r)�(�[q��Zɦ|g؋ر��=�<BlH�%:��3#��W��ݚf#��#�
^���	B)�tL������B�m�s�|R��Bn�4�"2�=�G����`J��';\N��j��G��|x��ac��C!yY���'�gR�(~�i�������@-Ӝ`�	'j|�J=:ҎH����0��\�D~ھ��o�z�m��jbp��$�L��abf �!����_�f�M� H�b�9{��vX� =��U��|�t�C�M3��_�3�����RI���-xo�q͉W����q}@r�2�05���2%��\I�A��k�R��HB��}+ 爢`���8�j��Q��]��$y<����F���X��a>�8~�0�Ϩ��f�qND��6Bc������L%��M�\�ZL|�4{_�e��&�-5�= :���Ӫ�T�mK�"��WH/lo��!�G�lif�����8'��~��J�w�i�uֻ�ȭ�Y�Q�� �0�p�;Z�Nf&� ������}˗�-��wo��0mUM�u�&ʯ��t; q�����Pg��s�Ja����J�}�T�0�)��̊�jf��w��Z[��Q����\\��żwt�e:}�&2�,溵��e��e�|]����Awd
<��麸� �K
�L;��u}���i���W?��$Q^�81���0�;~[��|W�4���c̏�l�ڹ(R�&�7e�إ����XQ!� �6��xZ�e$�!�����Ok��)��w ⟏-�t���j̐�h��n6�G����1���sHԯ�C�+�����]y.:�҇I�*0m�&��j��7�H��͊(ӥL8s8�/�%�]�(>��x�J����ڪ��Lڪnv�&��$ �R�XQ�zq�@%C,C>��������qCGC+L6����6�C� ��5.~޼�b�B��Q-�e�-I	��}H�߾S���B����2R�vt�RO���$O�
,+�*%�	���Dd�W�{�BS�K��2Ξ�(�e����JM�n�SS���d�'��x�/e��5����?�N,��b��"��o�QB� �h��NnT,�ѿՌ�o��I/l�s=O�5)$,v�I:��/QpF�cZW�x��=��?^˓yL�^__s�e~�;O0�u��)V�A��C��W�����D�2F�d���=��g�x�׭
ĉKpR#[d�O�h�1u�`#��N��f���Xz<A��J��W�*�,�	i�5VȱJ�hG|1���o�}Ü�c���Ac��t�7b��3�����O��b�,�½�c~��6��Ť<�@[�w<��mB� [�kqA�F�0���q�P�0�nu�����(֩k*ָ���y�J���I�Q!1Vy]V��7ciJ��o�0 f2���D.��Xcy�i��'F�0 8R���k�.&�ɵ�_���5Nי7���"�2��ȏfp@"g_��u�8�5a��p6H�7��ڸT��x�0�q��?MZ�w^�����Yg���C�����ww[W����c���A	�_�P�Z�z�<��'��P�i��,�в�o]�!��y��)X���x�.���X먥wa[��3
��GV�����S�ύ�mI�_����m�GS��ν����N��>��%���������hMu,";��Şrj���i�FMF���`�*���=�J�Y� K�qj�������T�������Or�kc�Lb��Us�:��N@0a���M%���N������@H9U�����ox�Z|�(B�n��3�	9�l������	8>2%����n %('�%. ͯ�S�݁����0n�`Ij�f�K]�k�V��æ�VD-��O��>�]zL8��G�ɴ��-#��BL7�/TND ��n'k���B�1�9��ᦷ@t5Я��M+u�����nـh��~h�9�����IZ��"c�1�5�[א���$���_P����%��q�y/��������*�A�Qv�=V8�B�����i�s��1�\��n�T�|J!BR'�t9;�a�S�� ͅ�H�H�Nߝ��g>�w<w5#�n?�¯N����Jخ�)6�v͔^Q�4��8Tt�Ox���DM]���K1��Ϸ������m��RS,5B*��|��Y��>�^��A��F@`+c�S�7+��-Uq����kC�DaaX��� ���
$�s��Bi[�4x��#j��X<'40U�|�>C4��c%eZ�#�<��7(��ZE`M�o0���Z�h��Yw߽We1��69�(l�ݴPC^#��&��)>�2���
>�&S���	шF��zD8�y����8�	d����5�p��v�#!\�r�Z�p�i���� k�A�5�Bd+�,,vu/ɤ�$դ�Q���0AӲ�ַzҌ�������DZ9��_F��e����$g������~�9!����� �0��`p���m��q�;��d��t��d_>���!��	T�;i��J���-��-g�ae	__A�"R��{<�)���0\\+I~u~R��,2�H1�A֣��PӤ[/�Db���Ag����b�7��������ȃO�u�~,��K��V����~�_y"oү�R������]�h'�ι��/�7�-��u�W#T��n+���Nv����h4|P۷5Q���B��M�.x�a~�&n�N����*��dN/���U�U[�ɵ�mDs���罡��)m��v��c����W�D��"�)�on�|�)Rst���Ď03I���#�FY��o��~]Bs�#�^2A�Ķ��p`�jL#p<f�.��ojS'�1�d2�",_�f��9�	T	��vE��5�Y*z�v;�*(UBj�瓴ǥ� q��x��1��$��j�Nމ>�RUrD=�$Q�_3eKB";p�%�U����
}Y��RH��۷3��t`U��}�d�i�3�e���/i��Iw��,6����#{m���B��t�5������	�:wD��\P��]R� -���Cub�t���BI��r�-�3���y+\<�D���0�����<�DZ�5!<Z]��t"��4C�v}����=&ɳ����ss/��c_�����_�T�y[9ÈN�	9�u�Npd�N�#Wx��i\IVd^���gP��(}���B�n�ہ�M�.����7 ����-]������u�٤�+`FU:Uo���RJ��<�����L�M���ef������z�3��P�� op���|����	���jE*j\��o�H�A�՜}]�:�����؍a��O��I���j|T���~Q�aݫ:e��%�P��:�)���ETo� ԅ�m*�{i}��%��{	�oBI"�h$���zAU��]"��'��|Y̪�ԇ���P:��'�Tf�f=�pՋ�E-���^�o�[o��;��┠�&��wři�"�8
L�1��GP��'	�m��1�~X�LY��X?GTf�)b�m��O�-,�i�����$�� �Ƨo��w�m=1�$��W uw@+��j��g!�()y��ԃP`X��{��'�e&P<�g=�iRq�D��d��K��-�K�X�(Zx�X�/%�����4`�
���������u�k��GH�]\r��dы��y;���^�(�+��{^Օ�Ii��80
u��*����ߌ�:��.�
bX��Sc��sޞ,l�����Zju2��Q2���	�J��D�z��f�Cī��N��4Nmgu�9���ʊk�6� �S���)^4�)�m�Y��`r}�GB�:=ȸC�>��
�U,?�~�h�9���@��h���5ҥ���&�#9-I�L��0��j�����ْw�ʋ�ji���w��S����#Y������5��k�Ʒ�0��,V����"Z��y9f=��U��7#�a*sYcCv�p�һ���VI�im�������P�LI��0?�� �~���g^?ō���i��Д'~�E��1R��(S�kH}1��*Bx�,T;�eY/�n�f�k��a�pj]�t�6��a�l�Z�Z.9�ׯ� ��>O5r$a_v�b]��AQ�kw/��e����*��("��ߺH���#��dwPB1�� $�9>u=�r�� �
+�\��H�o0� ��̽ǔ�����S)�%n���˸&�o?у�+���gY�t /��tR�i��j[Q��l2�EF�5�>
�F�;m�s���7��@IbǙ;�����L ��o5D��:�g*p�~�w���,c����;R��z�d��էZ��;�p�\�����G�<r��ۺQ��?u�k�0�i��.2R��t��
�QP��ST�WlG���@�,���^�?�ߖ$긶|�z��/i�o8q%;7�"����]y��k�vzG����:��F)`�n�b�O.�V`�Va�VJY>y�ո����[l�h,��9U��C��vт��]��{�N��!����}�+Hnd_D���y�7��(�mz�*�A�baw.L6	mC���y�mƿO���'+ڭu�Z��cX�U��n��>��.V՛s<��sV��!�`\��y�ƞ_�������;:bl�	V)vJF�����s���Pۈ�)/���S/�&��I��˱u)���R��k��ɾ�6���1�$)yV�ٵL^�9[SV\�M����zx>I�O������wgç��x�x�)�Zg�X��m�5�����Y��~=��ļ3�����[\�2���`�h�n11ƌ����/2'����|���/	�K�˲���@�\�'3z��,�� ͭ=?�I@�h�����dۦ�StVG�r��0��c��s>K�
>�~��r��k�F��Z�ܽ���B=�����`Kڇ��`��"t�j���D*go�[�o�Ɗ*�zL�K�Ժ@`�UXk�:_�f�@w]���Ps�Mnn5DSrt-�s��\���$�RO���.O��+�-�kд�R����D�'2�&���T�x�4�sr.B^kWA�ፗ�a�#)�~��I�'�A����G��̪��4��'��!P�K�B?v�t�2ݿ,\$.vY���#���Ӏ�e2�Z�7�y�����:�����*�Y�{⻓v�#ZW*uK�>űEE0p����E�ʹ�_��Z�XT}m��+_F�ZI����