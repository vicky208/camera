��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:�Q�z�n2�H�U��θ�����crH����;�$E���ê��
��G�W��
h[��Qd�+���T!��4,3��*����(� �g�",y�P�_���Ɔ����+�Hp -l���5$���"W���8ky��s'K���z�BD���0�gNr�Y�r�wre���ܑ�}&8�j�g]X	g�D��O�D�b=��+!I�=�X�4��&�����B�ε	5��f�}L�ϩ���=ɨс����u�\�Ȥm����t�H�/|bx��t;w��F�(FiI�~"0�+�fC5j`�yRd�˲)zq�D��iX���vH�q	i�wb�
��t�/M�?=��^c��"
/l�����e�zS3��u�KNU�a����j�w�_�ti1�<���ig���㎤"���k`�#�u�����,X��$棉�X�F�D,�uw=��y�}�]%1��k�0��@���9�+�i��@��6������d�����S{	�Jc�߶����L��u��If1\F/(�'-gy�Bs�X�]�¸���G哤�	�KhAUPOuy��dM���z�%OY0��/�W_�������D��/�bN�MϪ|[���h"�G�
�0��=�6�}��7�{�oKkʘ$
�:���_��r�⎨,֛���0�ǀ�t�.���4.�sz/YA�ì��D$�fl4e~<{ۓ	T�a�	:�.�B���~88Ÿ���,�*�ic�+7E"-�B�ئ��4��q"(B��f���t�.b1C�$K�6M�Qe� ]$�b#�4�yDjRq�#�+��- ���J�ܪ�Q�Ъr�I~v��b≕~�������GߙE�Z=�/�:J�_Q��MB_�dh'��ub���z��C�C�f��?�u0��у����Rkӯ4�ޫ��d޹��r�~&-)Q�7݁���a��!0��I��s��%���*�%Dj���	i�b�
��	.��)E.�9?����J���f��m�2��\�T�_�0Ə����q��u�&�h=� ,N���ps���śT�Mbg�Q�75�t�\q��u�X���_xB܌S�)u-w�G�����/M���f�1-dL@��3��;έ��*�OgM���K�1�3�}8�IHjD:��E��{��/[ 玬l�����v���	<�N51D�t/��s� �O'j �q��r�n�}pV�����C�H�x�����gR��G�~��kQm��۝�_�2m���W)y���5�J�t��J�P��W���;y�f�s^��sqʹ|~���KJC�Wl@W�����5�c��\�@1�I����x�����̇��f�`IJV�v�j�[�)�,��'}e�'��0�'�J�>�r
��CCZ��2�Q8߶�o���� =�� LY�sd�6�]�4�R�B��ԉ�� $���X&
@ �0��;��:�.e�Ŏȝ�(Nh�|7��� ����.v��<�����A�������d�̔t�"G���Z�y�$bR��y��H�C�q`6@�$eݫ@ ��o�����r�����r�
O� ퟵ��<���Ʀ��c(�B�UYq
O*2̔{�#/T��@Q�/%U!���D���j��t��.����I��������EԹXMp4�d2�{X�6&�/^�M��`ȝN}��#3��.���
T�JQ�$����XW�����}���T0������_������5�d�Ɗ����l�$���ah�)�o�����F�\�����~  ܉'�f��C��JY;L�\�	c���i�,������[�<�
Y�0�r)��i����ラ�v��I�T�a�e;i��^}�E3'��C���kN�^�)���kw���2n��^���-��}�Z�γ��la����r?23�p�P�5zk�&��~���@J����l�x�B	��;�8Z��AZ`"�o{���P�,�~&8�!FW5];CL�fZ��V���je�.���orTl�ȟa�o�Kϙ@G�)-b��� ,���|`�${��2��6=��0�S��	����U%�!X2��1��zHN���:���=PW���	�Z�Mv7�ڎ�$�s�OUh��ȵ6+��5���K/	�;̍7��a��l�)�wr�}�$6��]�_���H�;`V������H\T{�Z�eJ0����4K��x֪.BuR~0(c۫�u�b� �R�~.j�8��c��G"N���h�s�-�ٷA~©�F�l��0@��)�T�xO�r�l|�f��/�W8�t���Gֻ�V�~_�u��6��:�ă�:�Nj*~��4�{��y!'�����	��2�z=Tf_�D����w�"�AvZ	��������r�3��E��-8�-�z�E�*�"
�!%@,!�eϻ�Mf�͑H4��<�5*�~LBE�"�H��n���^���!�ڳ��S�4�%G��5s@jA���_B��0L�����}����ƹ�<��)�#]R�Zn�*ǈNN;������Iޓ)sywU9�y��D%�\H- k�UT���E�$"�!s����ŚMa-ծ�4W,b-� �qxA�00�g/�r�Ƭ�X
1�`4���5��Gt??�+��|�83t(K��Iu'�Mc�p�{��pD�e���w{J�&��P�{�H~��kc*��X�
�����D�@����,�B}�:a�^/5PO)!A���+�*B�
5��F��b�w�Y�inU�#e��/���%���b}�x�d^�~��h28W%4\�&|g��0���h)rm2_��:�B�-�D`��*�#�Nr��O�+�䰦��� ��`��ܣ�����}8�i4���/.�ڍ+��:B/�^���Pp�4ݽ�E��^\^;Þ7�D�3��l�4����v��|�aTɰ���8O����{w�'�7��sC����]�m���͵����Ŝ��wg#������c�P�lqVG�{ ���[�9	�ՋfԵ5�W6k��[�_�o�x���p�A��`��e+�D�7�UuB�Zs�����
%�0FzN�~}�/W�fk�/&X&���0�b��2{(X7�κ����v�Ҥ�(�:�O`M����[�q�y�gי�Y�����0�uSN��4��GB�uiR�=�)iWjE��oi�On�~���ha�q�&$*��L���'"��l�:�����Z�q,�krO��BT�I%�q�cd���<UH�O"$ь��io��6Fl���t��*%ޫd+���p��xG�����$8h�N��S$l�/���Ʃ
:�J�w��,;��%�)��e�n"<n���y.,�J�y�+�a�~x�'��-ϡA���~eZ0�(�F	u���MAw�{l�Jb ���*B��m�O���Ϻ!���2'"&�
E� �� ��s�yX�;��!_R�~�8�a��u�)��_ӈ��)����Ԁ��%��^8�c{M�����7
��i�j��� �.zTdw��J��f��?@͉��zE�swHjr""<�8((\��8!D�7� �2�CL})��n{#�Bį��2��hE�H�J��#uR���E���.:�k�R��N��N���~���Q����00��Q�e,�d�5�R��I=B�\�w�Y]�N�R�2������W%�cr�VG��5&|��,�w��G����u�#��4h��Z:N1��1���ר��7�}�/�ẁ���{��w�i��®,d&�'W4�!A�������W�1���8�;�m���q�����'�>U<���|�ɔƈJ>�	c��h�H TD<PU�q�z�	e#�"��i���G�I���ʗ/�!R�J4�(��9�ˍi��c54=X�͹D �2���K�u� �{�RT����]Q�[Qv�p�@s���<�SgЖc	R��촪^2]Gb���\��J߀Y����^��d�f�t�#|ģ�+"�����X1��5|H��T����)�����:v��Ә	��"�E#������|������JW�:��&�GS���]xS��Q������dc䞻e'�U���\����l:$)ܘҼ`{�^7P-;O�I��sv�I��'e����Q� ]�R��tƢh���#��;B��A��	5$��dXRVC��߯�&��~��Ș�u�(k�x�
*�K��=l�%G+�S�'p�V�Ŝ����{�0��>��T��;�-~y�l2���;��玝<�� �tY���Tj/������d�>�������V����Q��\&i�~���s0{P�_Ԟ�kj���e���\����m�y1�fx�k[dI)i��y�ζ��U{���%3-H�;?����;'����2ց>c&�Y&!��L�Qy��{s������N�?�C�1��(�����5�C��T��e	�j,����ۢm���c�;?�9j`��+./�X��͒��5���C.��C���(����\0��~ӆ��}���HQbYV���@_*b��,��tV��rEHx4�w�o��4X�IԐl�d��v��FSO����^��d=�N�=u�:_n�W-m��9���Ҁ{:}��,*�zY�v�����?�oh^ ]�YZ&�c�⎇8�C1��H�Z�~��MJ�%f�Q�?<��w���7��{P�ϥ��{�*IQ#����ԍ�ӆ���&|j��3��daC@S���B}����7����I�h["K�CQ�&����sS�7���W.�`�:r�;���8����!^Wb�^<�ݧ�,�b��d���U�yu��K9����n�-��{9����N��$�뗵��q�	.�����u�2ro蛺��!�4mҰ�v�ͭra���w9V�`�}�
~�ˑ�� =�Ԟy>.yp&�1��J�p$��� �H�Т@����p��Y0�9�7�RV���l�3@���_q(A�LC�hb(!���Hba��� I/t��Ռ�L ���U�{�>�@�X�u�-h��P@��Z�Y@��VjY`~�~�B�HO�Q�.��0���۲g*�wZ^b�$����b��*t1��k�����!�A�y�#8��4�0w�..kt�h�Ԍ�c�u�y����y0�fS��]�ɒ��rS�G,�=�����_@6سٺ�����̓���o���O֕.h�B"��*��F��J�$$HԊ�Xk8K�T=�q�.N��D���q��O���Br1�:d�\}�k��j<#\l3����2C#Jg���â��%yV�U�٪��V�3 ��U�T�X��N�nx�KIcTQI��X3Ѷ����i����.�m�eTh�L���q�hAn��T�4�PP�� `�u���cN�vxK���?r�x�He��.F�i�Ӏڗ�?�=T)h��t^l��1���S�x�;�1�s�'F����(�h��VJ�F�$�|���7$�:H��� O�0���Ϋ�`�}�I E��&�������z�by��-2����-��S��y.l��