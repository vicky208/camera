��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�U�v"�5���rLRU����{���8,�g�1*��)�����Vh�4���[*$�v��_Hn7��,=��R3O9��#��2@v��H�(Q����nQN�%�B�G��8y�6�m(˘H�KI,�K+5$�2���m��n1눐���`���1R^���A�f����b3��V��3K� �yK9�ܩ҄��E�a����4�2�{�Zo�x�mh��3d���<�� ��Э�A���Z@C�Uð�eo�5-I�+QZQ����9�v���4�0�l�!��[ 1�B�r�νs�;E������w�,!>�/qvc�ښ���^T�������~/r�Q�X{�ϒj�Z���X���y��n�1�pԮu܄Lu(�qc�`����S������n�zr��:e�ٝ����-ɳT0�,�����<H0;@Ɲ<����iٯB� ���4��X"�U�A�k㓂0T/�=>��`tbI�m䁋�Dk3)u�A�Ap�>�m�����1�rF�rr{�`�gև`}_W��f��X rW%���Փj�-b�I�V&���]�N�L+�"湋!�]�&ѐeX8���D�s��p&Q!7��m�*)>��^�:�����t"I��X@�?C)�(����dǉQ�������ʄd��)�ßk<;�<-;?[�ս��7¤t³�^����L2\Ӥg3�$��^i��.BY�p��w��/
tB�S�ԍ�*��"'�@���b�P�z�B�	0����/�@K)�zЈեR.��������i��[n�a�7g�w�c1�
���}X5����Pi��Ѡ\�Vpʐ}!xP�w��|6��Ӯ�Dh>fe���ۏ3�� K���<�*�����ixϗ�y>���i�F���I��'�YJg��Z�o��;g�:J�څ�!��_t�S�"x=�;q���}��@_��j������}`m�z0TlI��EK��^L�9�e �	tI��޻}��a��6I�����9��P��-2ius���}���8���<д܉T��e�$�'Gٝ�`�mS���C��о���/Ѿ�q��~��TZu^~�I�� �z�ј
G���.���\&:E	�z��&=��	�����-�݂G�NӼ�5OV����k�ȭ�~���>��b�G�w����_�1�"�E	����16i���5-�|��J�}Q���h�K"�95à����@X�"�	ޖ6�k�A*I7��B�j� ����i!ƟB�}ċ���9
<���5:}q@�-�{�#U�cW��/=ya��L4Xz-:��G)�ҁ�_^(�>�0���#�g,5�n�P!�y���1�V�r�Y�8~���\�7Q��G�)����Aˋ�6
�K�*�f�����s_���O��i�v�Aڌ�0�*S-F��5��8��+o'��y�� �E�����/p}Wo�HN�_�6Ʉ@H��"�5�P��W�]/�4�j�u��^rܣQ���UQ�ߕ�1T"i%$��b�H������Gq�2jӄ��G� �a��l�X���.1K���vZ��,�ЀŒcu��Â�
c�@H��z�΃�p����l�O�,�z���P��  ���"^h����w?."ӊ��h��zd��c��h�1��k��JD���w�pL4kd��'�C&��z�o�$�f&�l	`A>��]�NƱ?�ޙ�O���V�##�OL��ޥm�&��<��Y�5�[�͌L �q��τ�Ȉ(�%S �0o�Ô�ƻ�pu�'�~����v0S
�;���(i����h@�[���N�XUF�6pX���P�~%���G������{���g��{������¨��Z&��]��aE�K�R$��$ �u�Y%�M
����A54��yQ�K9kRl(�[��Co�㮔@&}E	�j�?���֋`�t��'�c!�1�F=�a�Lό7����65�h@�yf���-I-�_`՞��˽vk���IzYΧR�'��g<F�M��gQQ2���/��[K̴	��a�`�%┬O����f dk"+��~�+�xb�__j��T#��3|4Gj�^Z0�� �ZTZR�O��^`�Ia���S��܏7�ho"�N�1�@x�Lt�3��/��/����ף�b���c�ϓ͜��p=��������r��_�`tuZ����X��Hs���e�3�.u��K��S�I���y�ZV-)
��P�7j�������"7�'~�vT��Å���M
�������#�P{���s�ޚ"�z�������h�
�n���S^���`IU)�(�n� ���u0#~��Rt:9�4�����9t�wz������3l�E�1ؒ�Z�7����/Or�������荛���v&e��	r�jA�G�zs�z�(	z��>�+f��U�Wh�F���P���C��w�[/�qd����'/KB�����
K�@6��K��8&Ft����ڬ�I(�)��ݠ��>,��l�L
#W���&a�������$gj�m�J��O���u.H�H?�ص����W"'AϸE�V������O��~L�2����l� Z���iZ�q�zĽ���o6v+4O���{��X;�m�]	�p�]+��:�#�'�֪<x��^Ѫi���l��!K��4C� ��_l'��O痌ꍪe�y���N��RH����{��Ѹ�LJ.��1��):Ѵ�2�ً5f2e�x/�	Z?�l��"����1�TC�K`��d81u��Y�d^��GcـZ�Q5}�PDA��t�"1M�f ��$�3��Z����q�!��}�&���	�/��u/�>���߈�~h}��.�:m;�SU˞�p4ʏtX76����@�*�B�z ����z]U�?��
��1�h������
z���9Ϭs��لG��.Ӵk��䲴^����|&a�x!����8"|<E�� ���2":��b�XZ��v��!�3���&�E�;f�u2��@��i����?��'2��J�gm�jVU�KTd�c��p-�P��3��Ra�q�2�6�E��~��=�_�ɞ% 8U���L_1�xWV8�l����b��ɔm[���k�7��U��-z�E�����/��������@�&��M\G�5�&	�,�!O��WȲ��#,�H��FOۧoj�goNʖ� ����Rg$+�<�GP���;�>
]A �͢J���[�f?S�_��y �$�3�A��a����)v���3	t�+�� )c��ٶ(ޮS���=�	{������..hc���6���_���"����]�w.E|8Q|>���Ȓ9Ԍ�͓�쭖�l�>��l�Ҷc��&*oQΖt9�>6:�6 �V�2[�u]J�$��W�����I���	��Q�.��<ih8c����0��M��d� ��;������cM_��p
jF=��r �\���;���{���A�a�:����8 
1'}Ttz?׶������p�qƤ����e��#��f��Q�����j�x����	H��ݮ��j�*��V�����r}�,������wUQ�y�%��d;~Ļ��wܧr���[<��Jrå�E��c�+�����q���?��Ncǲ\��i��E�@����Ε_9P�V-�P���*Uѿ��-��V�N�0�»K�v�6����&��������2�����0��l�d�,�t��1q�j9�<�f�Z�y�C��=3fuR.���h\jf��6��I@�s.�s�iF�Y"��'�e����i�f�#o�U��4�r�&|Lt ��ǔđ�MO+��r�.����M���Z��&=2��9�<T����q'�����q`�ٹ�5���8AJ������%a��O�ʳ5�#�=&�Z��8Ƙ* r	���;�8c�iS=V<�7v��	��PMN��-�Ͳ�����+����f�re*�_�H��(�R،Ke���*x������bIA����\�;��		�R��46��h6 oqr�ye_�T'��(��5�Q�.T;uiK���b��z�I���T��o��(*`���zV[�S�GV�x�$us�V��"�'����4v���y
�hk���	,K��������K��Ư|6�+����Y�$�x��b/�0�Ԗf�wW�D�W��qh�ĕ���4�:~����Mɦ_qi� r�����c�D灓ף��R\���iƜl�����[��:��U��1.����.�Ї�9'*	��jp� ���FujH=D��&�_��
��CF��^��<����̻߷O�f%ܙF����Y���me��Ҩ���i�IE��k�;I�Z��~@�g1��H=�[��+D<p��oj��V�Hw��_�Y��f�b���`���~,uBwL�SG&����`���z���\�Q�nc#0�אCh��V�c�=�0| �/\�������=y!e�f�O8D�DK׬ѕ�Q<��2L�`ĥ��M��+���g�mk���4:�2S��^d���Zٹ�Ǥ`*�5��u%����a���֏ogC��:������U�8�-ִ@�p�U���-q�$�@�/>��~#A~��ɦ  �^�E��S􋘿E�(��F1�DB�t8��o��H�qe�ʊ���gK��V���ed�Ӡ_��H�a���?�<��%'�6�0����mJ��Va���<N�h�Pʜ�q�)��>�2�#�|%o@O���9�	0�"�X����k���j>m��琷%�*�zt�CZf�9�<=�2�%��HRǲ�	�1��A�Ljv���
9�eG݋��������`k�,Tr�`6�=A%�'G�c��k����P�X���'N�h]�ɒ�2ș Sڜ�X�:�l��P�Y[i1����K0~h2��z�`G�]���f�
Īs�������1 ��5��W����# O����������įb����p��te�z% b�	���Q�ЬӅ9�se�<�-d�2G%�$�:뚿(}=(��s��f/�ڙ�F52U�~_�;��uƥ��bV\ֱW���~��UUd�</�FW!��UI�X�V*��E�h��t�Y�Kz��1�f� 2/p�'�c��76���4���~b����#C �6c2��{������&JW�0;z]Km������n�3�X�p�qآO-��#��|gu��
�/Ϝ�&���_.�bn�,��ߦ�ma-K�ےG4��֝����e����
�>O��Sb�`����q#m�q_fz�F���cZm��a����~�g��/u8����w�g;jޅ~��E���nR
��
;;���斚��a.��{�M�ՠ�v7ߋX��CH+� �:��D�Z+A�'�y ��!��Ò�Php[}�j��T&i[TP�f�=1�o��UZ��>~��?��f�}�C#�Q�vlћ/���G��n�l�GDk���Y�C��2h�.�U�YÝ��`���U����������[�ǹ�
ń�lb��:��j&,sEd��9g��[����h �O$�����tƳ�)3�BO���s�vh��N�6�!�"��tS�����l[ �fh1}�O�ܨ�⡌��ʠ�5RS`M���+l�kj��7��&E�U>��������3p����%�/��,��5�r�`���wv��xA��&0UjN_��+Ӳ{No"���3;���Y֖^.4�p=��\���K���_iƤ�Θ�"AJ�⩁��Y�$<�|�1	��d3� �T�L���D0|�?j�"+�(d�%����s���4ɭ�{���B)4q-���6w��hpl.�;2G��\�7����I*���n�39snN@=�b#=�"��Q����*K��`��3�<��H��ȁ�Sc����Cq�ԑ���Gc�{��}$4p�Ϝ�f��h�����Lj�c��ɤ�έ@��y.2�=�n�`��6�C��/>΀紕�2!���9�Q�o8ƳM���A-+���,���+�����S���p����E��j{L6eF!���R�Y �> �oӏ����P�ׯ�x4���H�>�y=7��%`Q���5��!|ND������-�c)���;	�U�:�B2�D�N��pz{cf<�f֥@������K� �C�𑦋�S/�7$�n��ζ*�=�Jmy��K������6�#�6k��L��##�x�xA��>���B*ɓRA���Hk���U<'ˢ�}C���U�m)���_C���g(� ���	UA�>M���^;u��.��;;5dSSv�.�eE�M�2Fs�p�Y�I[X�d���S�[K-$|:��&�c4���ؒ���E�v�Ep���2�sb�5c���[:��,�~'ֳ �t�Z��-�� ��f�`�^N.+
u#�V���w�Z>4<n����������;�S%cW�����Hz��~�\^����\�ߏK4'�<!T�7� .8r���m��u `#����C�7Ⲛ���X8�[�g�w��a�p��/ ��W�_Τn�34).҇hs��/:�:��E��r��"�C	z�ei�g�'	��c�%@KT�u���F�*���!/��r
��bN~�&Ŧ�g����M{t�\�� 2��Lxʇ��� Ƥ�u�ɀW��ŭC�i4D�VҦĜtW�����L�4���������br�9P0a�*]�������( ��Q�]���I����C��ef�Ay����%x^HX�5\6?Oi����F��C�<{%�a�|��%�#DIX�7���wQBۀ�2����oyfѢR�,=�����]qa$5�ާ�A���s�m���Z�G����K:諧@F���'D�Ÿa��ig�uh�&��,R��8ȆU����K!������\�e���o-W�Y����{���I�b�U���.��z��~Ӟ�f���7^��#�]��;�<��P�&��( k������I�~ ޒ_u��k����'�~p�oa�u��c�#Y~bj;&��G�1��-��	������9J�q�L��ک�-cZvT�͜a<aA��U���f2���_\�����C*b�.'�N�֌��1ZB��4�>vBY�m�_xZ�4
5s9M�a������\ig�&zOh!q)�2Dq�V�,�5��g�R�Z�R����2��lB)����V�I��*�HG��gL���~?Z�@��j"$a~���c4D��]s�V:�.�R^,�?Jٯ��SG��3$J�J�X��ync���)P�����F4�#���X��:Z�7a|_Ͳ~J8[F��jg�X��Ѓqey1hT��$�2����q�s9�* �$�D�^�rڟ�cYDn�f�7%Kr��ȟ��f��C��J�v\p?h{�H+M���%/�"waE���Tfq>�^&}�	�3m*)�G�_�5:�Re@�gmS���yG��w�)��Q�טo������u��цͮ���.���\�G���x ^�Q��g� ���#���$a�qcB�(�z��H�@��,=t���,�<�ϲ�̗�D2|����_!�t���;M>2�;搊l�O��N>���=P3j�j�Nz{�����������Z��չ1@r�׈c)٦#@&Y�C� ����l������L��*,�Tr���Ι�JF�"(�01��֒���S�N��q�Y�#��I������qշ�@0�N�j����L�K��V�tt�� 'p6ȍ��5`�\�N�(=�)�_�Ie�)(/qoе������MO���G�΃u�NRD?�vAf/I
�;ǫ����2=m��q��nˌ�/��ڍ�= _"������t���.���Y.��xN��LA�9~��Y���?���2��a��U�S<$:M~�³	��+���~��xJATn��+��4#�w�@�G��s�WV��Δ�c��<vU��@�Y�T���KNO�=�|j~�?��T�U�.��7
Q[RAX44z�sn�w�X8���|o��@D�7C{H�[&�� ���<��1=�!�Ǟ��3*�+@��TT6P���ڣI������LcZ��?���h�#zT�m�:� 7Xٓu����v�/��od�臚�Q�I(��c
`�������	R��<��1���ےk�@�H�+Zr�گY����tZ�\�
��m3dT1����X�R�n������<����x���yp����oK�fJ�������Z!���<g<=�R"
��ݲ4���H��	��KZ��姌�k��S�9W3n�0a��BNG���""6W\4��X)�Y�0��l�s�W�`�����W'�����]&��6�~S���<�v����<:��0���k�>�}��7���틙��.E�R��ˋ0�vE���|�YTI`�"�"�{�U����{��MJ���4����~h������~��g��J�>�ɰ�g�ήg�i[��q�A��i��2�<�ݴ��&Q7y��e���c����}p��HV^{ ��sw��7$�9n�<���-���E$ߩ��b�����*mH��U��:��|Qn�A�n��!����(��D�`uߏ����) ��~���9�gtO�����q&6�P��8h@h9�����T�t��G�R���4�wF�dVCs�*��p�/BG��'�R,�G�d�>�0�O᥹�Wi��_�j�ca8J�,/��~�3����Fz	�X[}��
@��J�t��b��j8�d�xc{KO1�Z�!M���Pm�M��fO���ptF�~w��>�U)��Ε|2���5ͬH�o��$���'��_��>�^���[$[S��n�����g�>���G5:�˅:7��&�b�ʅ&CT׹�բ`��MS�������{���(x'�������o��`�o��p4���6�B�M@�����blN��c��KT�g�����̲H$"�X+5{�`�2t�E��(`�X�=���I6�k$���^��o���߱2���u���
�%���^ٵ~?��Qz5X��MW��g��5ʒ��U����C��opM0���@.�$�'2=��ZJ�
��e�G��̐Uv��ңj��k��Y��ӹ�GD˕E8���F_���7�𱤐��u&e�*��ti�w��>&&�6x�(?�I�!Ю�pgҿ� E�Ċj__��[�A[O�U֔J�Ň�V��W�)�-�[O��xp�D!���D���C��k�8v�GbKI^x�k����}���=����c�B�M!A��Ʒ����1[}�{��pؤXX����2Ap��R�I�Zv=~��׹�>��jV�B���v�����_t�0�<cW~Ɓ�4�7���]�H(����<(<��E�n�iQq?��d^�z�o��!���+�t{��[���RľE���d�1��9��O]W������QL�-��Nso���1f�Y/�_!G���8-���O��j)Ղڟ����X��_o�/&3�PA��Λ�� �as�K��?/XXN!" �!l���+6\��<Of�����V��S��� ���)=�E��:CT8��00�Jzy����#��b�㲫V�������;�{Ai�BC��cx���`�+t3[ ��*�Lީam����@�v�&������l�7�i�H�+徰 u,���Q	Z0[*6T���J�o�K�(~i?�f7�O5�	��:+���:���q�e�-z�_��½YԵ԰������i��H�E�b�&nݬ9(T!ռ_�ȩ��>��7�Vu\�T(���<�2�T1�H_C�\�;��d�?�����-�S�լ���"�dP������t}3��u�>#��7l��h��y��ڌS��#�8��=2
����
��c�͙"E��w�Y���Y�@�EL���z\ɪ��g�k��M�t7�O��@�|%�ϻ��Å���a7�HE�pK�?�`�39�p�x���o�"��Nn� ���n��5R�LM:��t�K�}��M+����)s�yU�ǟT�&�ؾ��jo�#��`,?3}FF�Zk�©*�BhZ~h��/��0C���10�����6�vt���bC
�i���ȇנ�ԍ�om>Rs
��|*$���dy5MU����źX���ɬ�+�%��o�p��$lp���Yz\�Y��~�ٻ�Mq�#='R��@�$U��!1�� �:��Z�����RZ���&k1h���8lM�w*�ʈ������|X��JS��S@l֜.�e�5��hܶ;�z�o�>da"NT�%WT�5�������.�1g��t�^G4�$�C��'i`ؖ���]a������"��ꑠ'[��&jZg�ٓ1=�W�*_nf+��C ���r�uW����@?.0wro�J|=�H�m3���I� #�-[ΰ4��� ��`l�Ú���#S��C�|8u[��?>tL����\�xv�0V��q��|� ��v�~C��N�$���3��� %� ��ī	��v&ٿ�߉{�]^k���
�`��Gi���֓�*+F�-�#PmKkX�S�<��%(��_�ze��e���h�� ���g����1��k�����CV��%{Q�\��f�@:�}�'�B�T|Rw��MEq�ķp&#��(���ϛRX��t��V�%���>�x�4C�� �"Î���rt��V
D��d�������0��1M���{��B�JH���_<�{A
�;u5�'l.�˲�H�^�h�����W���ш	#�JO*V�x
�Ѡ������`�v���v��#sJ�,��}_�&���M�4����]�u�#�H>�=�4����|Ŏ-irn��BScь�r��O�Q1bY�.ل�n��(ς�q_�b��)�l%L|�q��W�졢vZhJ�@��4_Xe��Vq��542���r]%��B�*���^��[�e�bw�#�f��y�OCq�Wgr�|@t�j�a��ƯѠ�����j7~�<�Y	}M)k8��3���Vf5����˖aއё�e��o�7
�6F�M���Md1>���M_�T�KeՉF�D������\4��z��QW��*0�!	 �|���>�$��]E�s�͑TÔ���[bs�EX�(�t���yo߰����=����uvS%d�Z�WQ�B4�zEӌC���X��W�l�<�)̅�fi�W�*|�Ķ�qc�l�R�ٜ�N4�Q�����e���ǈ�<��'w�[Bxq�؍�&'O�#2t���6��>��&�{Y�FR��	�b'��50�V`X�V7FǖUD��扂W�?E�N� ����P�T����W�ԫ��!t�LZ�tl���ДOL��	]B����cA*1���r��hc���эp(+ƨ7X�C��Fu��pK��k�Sgߑ;���uG�*�a�
�H��F���	�>�٤4LD&p�����lf)n�[�q�����\�AN��D�l�XC	mvF�h��w(���!-c���؁�i��m����U������A=.����2��]	�V�Oq4	�晸y�OV�k�eU�݂ucj�C
F���G/^ЊP�]�	|A�-�"��^%T��]������P��9�T1,a�|��Q>�༔G�˖��ˏ5���` ����o'�qؗb�~-&�զ�ׇI��I6F����9�v�<����Ë���^4�80���N4�Ru͍�E>�'Eć$&����~l�*�1�]4:�`zdó9��!b%a��t���L$�a�a��T�,��'��	��Y2�a�T���m�n�&~�o�W��?�L�2n2�F���PZHUG�~��~�F0���Q{U�.���m9�H��ưu�DrN�@c���̔�X��p���ϕ,Y����`�"n�qB�����>;W�)5��s�6[8U^��9�x������J��!�!��W��%�]�=a����Mx1'�T��S���<>�nX�ֆ�NY��N 
H��D�����e&���ް���qU�!x�N '�-~��xhd��4,�} ro޹�C�t����m���'(/�Leܤ��s�>�{����ǫxG��S>�5A�ɯ���"I?����υ���X��^�R }�v0�j�F4P�a�����64���F+*O�ͯ!}�/�&.K�Z+VC�P*�y-�tU�q��0&��k�]?=u㛶(QSF��M���Ws��26��r�sG ��ZՖ�~PBװ���*	E
 &l�p�L%HB\��~�Ϲ�j4�}�G�k�
�34O@�Q��PyZ��wncR�'���(������~D'F��:���v�$-=*�ܹ��D�2u��0H�Ľ��9W�91��q9�&� �� /;�?_^�6VP(���6܅��A�F�����������"�ܢ�7^��ͼ[[ن��z[���}�ݓN��y`����v
6�H�`��2��!SA�����(7�����lc���� �QO
��I������Q*���OմeC@��eM�����sVN/(9�iγy�Ѵ��q=Lڇ�؈U�ҘmG�����z�k���&�}��N���d���q�hn�F���r�	'�p+��'(,�Ed�T����S��#���cIO 6����$T��V${��)h�J�s�K@�>�����J���C �aG���S��c�e�zf����� ��p{Gc��aqN8Z��T0����Z='7Mgr0�����@`�F��m�"�sG�����x��25�Y��a��՗%
�ݍ���e:i�~"g��a""��!eC�cy�[x���m�-� ��w�Y'�W�\9�����V��|�1c�����R�ジ��i1�wH�����}°�Žp�S��l:����<Zb� �3�
�"����d�x:�s�86�	׎J��V̋N�/���-�(8���3��6D���"D���nn[GY�%�
}�/�*	�ێɹkp�)�S����-"�p�@(�p�u���%�N��`=H�-M�|H���74i�3BԮQ��O�_w���B�>p|�Hs�B���NzN�	�qRݺ�8���@ESa�f��6J3[�[q�� ����q�f�Q�g��мź�2r���a���ۈ�r���`��ج�ąWxaJ�#���y&��d�zp%��~=���F kX��ddu�nO���9�!ax+iN�����
&�m]�+S���7���6'�}
��BmZ$}5��;���ˊ���y��x�p
V49��:H<���S3�l�B�@s%�"��ҥ��7d�W(��oĀ�8PHu��~���GO}-_j��TZ�G08�W '�3j�\��3V�`T~WɇKj�Y�nбܠ�[[ ~V�}�~	�;Z�cG�]Q���du�M qT�ΫD�)ܨ��Tl�e�^�Lm�z�x�rcWtB���<y�����0I����-}r�:��'C�?�.�q�V���i��۞ў�3a�!$ؑ+���7�9'z���El�m?� ���V���e��H3���H&>tB#S_7=ظ��E�a*�L+EARz��4"������C�3�Pq�ǂ�Z�flZ���r:�@��g$B�}��C�*�;�D��ܣP0ek��<ud�̔l/߿��,���@)�?k���6�d}S�-�&������7�B5����)^����Q�Fĺ�@��~�y�ƶT~^�ͯP�5��4M��Pr�t���"9@�*����Zv4N�sU�J�k��Ћ�C���D��+�Bk���L�2����`��q�Q�[t�j����k��-X{��d�_}��)�W�xj�x�L�0�;�{���i��k�����Jqy�w<W��0h�@���i���9�~�PXb��%St��X��K�1�� ǚٹ�j{�#�]j+xf�r��hΠ�)����;��##��B�&bըD�/Ͳ��0�|6�a6��'Ê�`g>:�#��O)����"_c�u�`'­&E�w�q�Z���\f�:��j���0	�
���8c���k�5�����C�)K�d�[��͗����^/G�*���Z���N�����qВ���ly0T��|F����B\M�+b4Hѿ��gg(��9�����rv�����x�
�>����.נ�ٝ$u�WK�tyׂ,�l��mj�O��',uL+|Y@���%S�&F#*]�S�O8��O�$��8�5��A(�_��Hl��?���I>�+�V�Ȋ�Y�z�����3��Ee4����G;��,���~�R�6JGS�9��@=�?�� K���'y���g���saB0^�-V]�����0K���\��� �-��$� N0���+��ŀؕĲ�͇zyYX�E���4�#!��7dg�H\3AZ�5`�Lb�$m���B�\n�'�K�)y�G��fg"]|���������}NtO��:`��.�{��ZxI?��c�>T�af>
�Rw!�_X��p�3��M�H�,Gߎ�I�i���$�B֍l�!)9Z%���B�Ҧi(o7?,ȼNT���A6(L���M}I(GQ��9��jlů{Zq���.�8��-��*Zxݘp�=���/��Q�����o�^	�](U��9������x&1��pB� B�ا�@�8��O8��P�$��T5LǶ3��=��Phq��Wz�@��$1Ew��4�u��-�߈S��{U����;�(9A�n;K�j	OQ��8W�_���:fIw\UN�u&�?�Z��U�\���~�Z�q�p���w�cڮ��lCd��%7}K��ln*0ag͘��ӕN���a���J�I
��ؙNڢ��d̉��D,|�#и�Ȃ�H�r�<���G粣q�Gi.io�"�O����Ml`���fWw&�Y>���j�\O��jaĲ�[�/ck�^x~Mʆf�v[������6��Ż$Yq︹dc�,��XE�uhD��.��N3
�nbc���*�8b��~t���k�~D�W�լ�}�Mʴ0���1��ԏ�R0�Wz�9�<o�J^!��U��4q���	�z!���S�Q���쇾#�2�N-��uNHc�:���\s��<�k`q�;p�6̺:�Z����-:�$��k���V_)�u��.��<2�*"/��ud�jr:+���� ��1��F/�x�Tb~�tё��6�Xn�5@
�Q̾w��9k��?<=�qTq)�l�A�%'����7ь�3
�$��P;���3��m�Q��okvu��T��S��ӻH��(3��v�ʜZAp�M%�AN�ʺ7�".��C"L������ru�	�"��=s���v-F�8`"�>�2Ȇ%�ѧ!��e .�J.�J��������������t�B%��o�H���[���P_l�7�V�2�%�^�"~"���h����;l۳j4�Cl�,�j{��#BM�n7x=��-��N�=�Z[QZ�K ��F���[�����I����U�RjT�˝�Ri��3kG�Ti�y�k��(���Wyq�Y!��|8�,�m�ʎs�~L�LLR�3Ċ��N:�ޡ8C�4>C����G�1�&�C���@R�'��@��>�q��H]BJn����H��zڨg�:��pH��Uc7I�"�P��_s�����D�+,H'�{���5N�K���[�\Tf���D~9�\kdxM�Cqߨ["i�uu�����PZ�] �O���y�u�k1&�QB2�V$:@�9�FJU�����������8 r
��v�3�*	I��`��c���9_2E�M�ܭ��ޖ��a��U��k����h�ݲ�"z��Ї��o�o)�`����l��9����,_���;�����?k/I�!�W��q9ﾊD�^�6�T>�2p�,!MR��#V�:I��Γ�] �*#vމJ;��	�Sg��b2�b��R{���4_R��]���"���o��H�Ҟp��A�I�n��_g��?��z���O��W�鋍rt| �� �DZV��a=[�Q�3m��Ђ�a?��T�ѓQ��}�RG#y+t!�q3?$?2�3=��*dW &�Z�dd�h-�=�D��_64�&�%,��;��I����*3Z�]��<{X?����K��a�."�%�h�
�(#:��WQ�&��P��p�}88�#fV�Pa9,�dƻQ4���RiTpH&�
���Spo��T�@�$��K��_,��瓙$P˔��',�M\Q-��]���aɊ�%R<��:��z,��FQ�St�����_����[z(pN\A`YbK��Ldx@�!�Wa���@7��%���Ɨg==��ezڹ� ��ө�^��kn�� ��Ͽ�<�[tb�%9��0��A�?Z�RO��	86����N�����2����T�Z��A+�4rj�&�q�-�r�,��7p��V���̥�:��<GG+��Y <Iwo!Yb�Lu��� ��e��k�����դ�"&�[O�ggc�� c���'n����Mѭ1���⪪^O�І�2�oh�UW\@Ƒّ$۰Єw�h�A0�C;��n�L��
�p^��5,��6a�ѭ]���H���t˔���-M�i��A1�M�=��U욝�Ęw�'�2��v�h��#TÉ���Z��u̢�c���H򞕊S��Q���畟g߲C ]������9��\��h��R�\`��;��d9K�A����QW�!
^���L�$};b���/��G4���a�������Jy�ʟ�CwuX��E�y�>nU�YHp3�]�&S!)篶����7��ھ!�׮J�r�ܶ��\�O�����逞K����R6w����W�	�M�/�~�5,�h��g�H��1?V/8�N4G�C��a�����w�����W2vh�"^��q㮪S@1�_�W����g��+��'����y[Ml�[c�*s���Η���1��.�ԛߎ��e��b���ۇe6	[�*m�-���WM��=�>�@\�O�=�M�? ���j+�Tk-��~Ҭ�FH}��$�eS���;#�s�.3�ݐ����[���ޓ8��4'��J���\#4R�G��wH�bŤ�� v��"R�0#�"��gB��t������|{[��/�0�}EX1�nKw[�*�
�����5]����vH��~=�(�X����Uk��	B��!v^��G�M��;�ƪ�kv���ah��Py��W`Q��x��f�Izg�"�����]��h�8PY��x+�\����+�=��Lʁmh,:��4�p���Q�y��k�%�j%�����Zm�!|�*���f��}��-Y� ��u��h�@.!�$7� ���Z/ݐG���--�[#�	�+5�oO�=���7/.b;Ы�2�2�f���s��rF(�k����X�/{��{�b<N
�nP{�I�� /���i�q�"{����v%��f 8��o�a���Nq��F-�Q��QK�u����*�<Ho����Ǡ3,�7���)Ы��P�mdz����Q;��|�V��1fs٭��E:tW�n���8kS%��^�;틢�� �W���O&�������-��FSZW��f��'��K�D����Ǟ��Ѕ2^rn_[�v��+dl4���-��简zGHG��H1�Q"|����-	Y����_�[U@����C��-
+Q���"u��?t���^��JΙ>]��Y,�z�d�R���fß��a!�쀳�)��_�z������H*��Z̧�A�N���-l�7���ۍ1���
� E?���k�B�!!ԏ�8�h��������HcS3�I3
"BA"����ꬄ���u?I����x�7��F�*�A��N���L�i�ʅ|9�%��I@ЁFR�؂���j�$ʗ�P��H��[;�2�t��A{�*�\\5G�Sl !Hz�<'��]�9��Vcp}�"���@����J�gY��|$����E�aW��z�+�_� �&�YX��{�$_	c)J	D���m�!�&���[�"�]35�z�n���4	I��v"\�:����u��Ѩ�j!�Y�|�0}f����bS�O��_
�Յ�r*��� ߾�lED��ts�ܯ�QX���!̠>-�u���Q�#� �C�$4�a��:C���~��� 8�i� �jB�>��J�л\�*�b���̛^,3�D��;�Θf��]1�YN;�:�_p��1JK�|��=:vwE/FFzD��>�q���?okM�13�ܗ"����n�)�V[�}CI�.䭬?�#_ y���`2L�팒�p�}We��X�".�CN���Mʆ�}p��-(_}J>�d�+�%��tu(��p�Ƥ�w���Xsblw�u��������D�/�ڟ 9�Ó#$ь��[v�ݐ���f����)��+�}�w֕݅2���_7.^��9��3~Q@�b�N�����T�o(��^;���oZ�v+���S�Bf� ���i6v�p��\Y�;U��bG�U���wυ�%kPg�BJ���:!C�]�Q��V�k�H9��C4��b��G��*�=8�� ���,<06[���LuL}J2�y,�`ro�ӫ���"�a�"�ِ�5��Hk� ��;6�kT��g�Iq�F�-��h��)���s?n�S���o�,��(ۣ���D��?O�"8U�p|C�9[$��I6�2�D�B�Cuo�oa�zI9�SB ��O�~�q�u~��V��?S4f#IA,|�o��+iO��O��e�}����zj�
��Vt~�f�:i�r�w}�����_d�Ks��<���p�H��).�9(c�IH rD��a��ғ�ʣ�¾���xN��N��fa��頦�a�.* ��*�l�S)��T�g���Bt�)Jɳǡ���O���W��fO�d�!Uń�?�ߞ�4=�U`OĐ�o��&����%u�S�,�F��
u�$@��3҄Z�% �WF���� #V@Bt�F.l[� ���^R> �M3� kF��#��~,��g���s�i;S�az7	��$&�q�p	KW�=��ߪ�2c�mQ���Tb��"�!���]}	�����P�f=��#|[3.r�e��-'1Q(�8P�]P�'�\�.��¡�,�OE��B�: �ڲ��=8���D	[y���r�7M�eՐ���u�.ej��&ecA�
�ǘ.E���{�!���\�|A�����e	�zs���>p8~uVQQh�������ak���r��Y:�B �Tý)4�I�,?$[��(�"��#��oQ��(ݷ��)S<���	�j�ĭ8�<^wo��2��p�l��	��5�_ۮ�l8��"�C���u��o���IH~��ML���Sކ�����L *n!���' �&>p�H�˟��<[��mG���%�9䖮r`��A�~������9)6���0c&�J�5����9Q}ی��NZ�TB9�Ç�+�u&����5a�t�����h�l��'/G�Lm��r*��[�oC �8*�Q�M	]f�g��.ė��=�?t#�p�!p��}��Z��:��]�kY�~�>(��t�'�\���S�Z�� 7�]�I������^V��h���̀�W�� .��t�	1�2���C�I�E08L4���δ�>۩������.��NK��bZ.`�WP��m�8��*H��T�4Cj����`���]���¢� 8��%CkzF-\���)|��_ku����T�6�U��
��� p����-;��2A;�$O|Y�̾����w�t̭�i s�Y�~�Hobl�_��u�i՜s
��P]��A�X{�ה�n4�HT�;B_p?b�k��Sa���ѥ57�w�5�ۍRN��ώ��1�k2�a�u/A�br���g�d�E��g<ྃ�A+�(��?妴Am{PP�� ��5��s$h��4�j�U�֗+����8K,[Q��N���(P���Ǵ��C��im�?y�|��eE������2YE|�㍻	k�����oA{r�Ɛ�p-�/��D;j��y��|���2����ά-���):�J��3ߚ3�8�&�;�TȽ��7P66���U��pU4�J.��|t��t9͡V�z����=��6rA6�y��jC�Ś��� U}��:tjRF�nx�g�M�f}׆٦�Y�p�l���F@�JK�mX�\�A,Y���/6JjS� ���축�eߓ)$��8sw^^��S�d@�Ckdw]�*�J�2ٛ��,�&U>h�0U�a�'��r�wnݚJ#e��3El���C
HtD�ȹ��8��I�:�%�l�K�|�]�>�R���]��9ӯ����p�.�{����T�|גs�<T��u���o���[�KX���3�"�/�D�O��i��k2�;I�[�cٗ��qU���V~x|��U��q@_�+�?�KD��ܓw+�BC�4���B�z�R� ����u[x�D�=�
T,����7�%�u5�Gp�^f�i0-~�9+�' �Q��6�SF7��ED�%��:�!J�8�@�����#�gNR�K
������NgY�y� ^��p�Y)�CޖL�I���>G֓����I[*B(5~��C��;�iǢ��қ�x���e�{c���l�I���O������x C� ~u����̢�k
�Y�����q�=#dq�?��'p��Gv��6$��T>ȱU��@5X������+Ϸ�{���k2�G50$"�%�#Ǹ�Ī�;�����d��`:��φ�ڇ�[�aLT���iA��:U��6����P�H�x�蝊@�]=csr�Tݢm�w��!��l:��]�v����Q��H������|�����a��ϯ�o����O��9yz�eW$���ϟ�8if-.�,�D{�d��)�ʦ���`���4�⬬����h)�����\��6�Z���|e. �Hʗ=r �=K�|�H�T瀨Է���=��n�1�'#��H�d"d����֏�I�������\̽[��$2_�|;~	�x�D���r�5�m �t���
��P�ј�Mo�l���dsL0�����O���ȭ2ٞR^ͮ������6����B�f9��������N��g��0b��^��Cx�KȺ�j�����¥u�<9J�0�hu_�R݅;�s$���6b��G(���IX���	�ɘGó���vż-�i�����a��������^p�@�os�/ѣ�D�}�Q!L;�����'�VTbNl_/@X|)�ET��3�����*0^a!B�]������L����w/z��C5*h�7w����(#1�zHl�85����*H=�q���Q���.���E��[ �e�6��E˂2E��9�Np.��mQ��tyz ��W��T^΀����뻧v�?x���s@lmbiV�Ͷ�Ck����QO�T�	͑�� �o�a�D������d�A:$D-`�>ݖ�*���&Z���	���v�Ss��>ܦ-MGp�|�[���p��t�̷7u�s�_0��S�3��)�}�W�c�H����A��������%�N�+�*�i���w�5�������F���5���1��Ag��w u6,r�BA��^����kx���e�����}�ׄ�2�H쭒��^A���&�'�/w�)�j�F�^���bh<��Pl��-��5��pTv3@>���2w X�
�\�x ��֍��± S`de�4"��*C��/�ȖA���!ZӢD�5g	?�~[=mnz D��[�ǨѢ{��+%ƹ�Lu��CU{��n�0&� ;�S��~I�ܑ�	�����F���M��y7f e���h)��q�e�޹���E8�9���$?��v��5�@���-�����dS�;<g&�5��W[e�Pf+� �֫f��a��H͟�4H�`�&���=��}���1��e�T��[H�>�A�{iJ�X�hC>�ZE ��",��P��s^�rG��Bf.'B.[��!U ���Q�%Zp'�[�m3�5��t�R�
�'/��A�����5�����T<��!��H���w����f�y-�ˀ� ���b�4���M� O�=qA����c�,�'/e�Tjq���XH�Sv���5�x��1��s/2%�\� bPH��}}����=���4�О�@�M��$韖����t%D+�92v��{�}�2���D^Eq��ի(���+��IPL���>T� ����?PB�S��V�(:ΪG�S�D�1\�/
+X���I�L�YD��2��eL�>ϕ���.��E��y�m������=)�݇���+.�a�S�F]���h���SQ,�����"�\ٳ��ϕ�tLnF�p�+0�Np	t�>u@Ը����L�* ����%���.�*����D�@�eR5�l]Zu�H1���6��,��4G�b�X5��N�PvtH�nc���1EI~�l����z6���Ƣ�]#7��[�
P8�৤AvF*e���z���
�H�@%�N����Ex�BkFי�M��g���g�R�i7;Z�Z}'�FD��ð��{(�!\l���PYi��u-�*L�=��ے��r�lz�2H�k�"�AI_�C��k}z�z�bh�!s�5��zC2z�����)f�������>F�`��r��)N�%*D8D8!��NE���-��X��F��p��}=V����ҕVj�?�ab�K�ϵԙ9�n�v�*��)���4G�u��A�)��cv#�~�����>�8.�@-W���Y����5�i�L&����`;��3�2���� ��#�!*�]�Ѥ!<\Xv�L����r4=�^� ��*$Ե�Do��fk�"T/44��s*�E�P<�y.}#�uP�*/dm�J?�"	"yw�`e�^�a�oK��)��]����N˺��S��m>� ��Wd�}R?v�f8��Lko��ii��v(6�Iϥ���yV�X��xh��+j�:t)�_��P)��'�Z�n�T]D�fq�T2ب_do�0���y���8�����ܝE��0��;���	c���E��HÖ����Zb&\����\�|F�̻�t���	,���U�7$�����;}��J�p*y�_��G�l���'f��ۀY�^�������Invx gc]q*x���"G&Z:���/���∴h����n������ï#e�:dWΌD�!�_���vHа����s.��a�O�B�f�h�D��ľ�E]h�������Ϊ|q�I�0i���bRNo~�Gĸ�i��%_�ӟ��)���9����b�>��	�)��^��}G�g��<.[��xqޠTQ�W�G$K����)HN��vʏ�'aV��QD治�au4��Z���(��V���,��������-��
������CS�]JFxX��~-�؅�Bۧtʥx�i�/<�/�'�scv�Ԫ?��5֭�C��P�4&䀨�r���q9�eVSڣ�C�Z����b�WuĬ����&��Q����f�[ё�g�Du�J��x�K*��g��U�;uV�̦��g8�r���� :��,B�0�w���}����߆��άO��I��Ga8�c���"�u�#Y�`�ϡ)���i����e܇���<��&��7�V��q�/q�e�㖚�j�y����Z^����X��b�{0��Z�jU����~�B�҂�*xO�}{L���}0�����ދS�?`��D�{�o��Pg�˞�ԢAU�`:|��n�~��Ԭ{��mF���ȵ�q]~�3��Nl�_�dYծ�h�A�pE�O��MC�w7�J�h��6B2�A���;_�~�E�{�ھU��ⵑ}�l_���3�ٺ&�� c�{Wb3n�g��QzOE菫�\�6VQ�]e�g��1��=J�a ���yd�Ȱ���dT��?�L`~@��^�	��b@D��;O0D%��]s� �͜~���x��Z��zu�w���B��v3���
��B�5��8��s�e���0�+ܢ�Z�pR'�tjo$��B��7scq��NªOb�f�*qv�3@���v�מ�59>V<���WA)އ)���n1~a�4�5��2-'�n���]���n�5�i��]�ą_t��<5nq�UnMK=b�^�����f�dw���Sɚ�#�3.%A'DU�3r�w-E	�GLK��#d��w_�|؜Lk���x�;J��<��%��#���{�$H�|�Q�7��N�_�t��I`5'�h����2�,�<О��1^�
��E-��EFjf>&CT��{n�E	�Ǳ�AM�:Z�ߨ�K ��~����7{c�X-��R������:��i����fCW��TK-BWDGGJ#��k���I�.�úH+W/��n�|\�Z���g8s��{G��D>@�����gs��͊�Y��d_��ղ��+<�����2��t�oY�L���G=�<D�=W���6��ybg����Y>��l��pkh|�����g���)����c}�d��&C�^�l�>~�`V�7�xė�L	�;�x�Q��J3���L���O/:zΛ����Â��K�ͼ��� N���N5� ��d����'"����s߇���Ă�;��]Y�"�{RR��U�Y�"�zy�zB�J�4φp�4񣎝���tt�����m���M�6[��p�u�[6�z�E��jIm&LN�'�[T�+;�����Ge��kՀ���u��Ll�2��PĦ��J��n�j�-��"�����2x�M�W��W���ٟHb���DFmI��'��a8�a�c��f����ؓ`��˾�3�v��ۜjĻv����9iC���%��	Crp�v$z�D-�%u�𨞛A	@$�J����&����*Z�����CD���,Ê��P��eԓ^iF�6�e�_����DW��7�$2GhzY���_���c6�B����m�9_�#�-y�!�u��(A>)��ZΡO�D[A�r r?����m�S�J���,uY2�b��r;b���2ZxД���X��t0�`����wL.���7T$}�Rj�=�̌J�?��L,�n�|a8��iw?,�绤�͇���/FE���c�:�H����?�Tӂm]��3�`.1H�@#�RNH7�b�Y�-a
봫^����h��i��Ʃ�U'�`D�>�?����u�y[fwZ��~1���HxRt�W�ްrU�P��|F��$X�ix�?��P��oB�<8��4G[�����#�̱)`�翇��o {�	+h�Z���i�e�qe��b*�L�U�;�����-N��JY8	N���'!u��h!c�)r�����b�ӱ }������'�V�d*���U)��1���X�YV̚�k�v�$(B�ܬ˫�:��e9g����֔ȲЂm��� ȕ ��Zy/�G�o�4>h�c�H��hh���]}��r�5�cM�9�+G�-�/�M��©���Ĥ�@��0��`����ས`�*~�d�%T�`ߙš�qٖFw"��Ɏ+��"�FZt�1Rg��=��ac��t�W�YL�@lu4Ċ���g4E����`�`T>`Bk!� �b��x�QG�?3���f�%!��e�Lޏ�����o|�j�]���T��`�_�·�&�b{٪{�4�]H�������hw:�ena�:n75������%]@?%�l���?�k�_�<M���׋�@%\Hq|rэ'
A�p�X�HSc�����C��x���K��V���
�نm#p狸�v%��·얌�|�D���ڈ�&i1��#�F�Nէ�\�KڋO�Ia�NQ��{5;`L��9-���iL�z�@����u�͋൝�fz����C7������uY�g��T/xV�M)�A���;ҍ��25�{ނ�ys!�Zw>]��A��K��Ɲ 3���{�k�$y��*U������3`LݫsÖ`='
FU̷��8ӈ�V4�/:�Um�������?T=�*X�G-H�US�X��!( ��?Q?13�a��ѭ�8H,Mkmx���[�EB� ��Y�]4"C�$&�lw��;6�i8;���������'�FS��=x��*t��a�����.uc {Į�����3�O8����YG�D�����T}߱�H��;�T���1�������K��s���v���i��'a�-8�k,~�3ἓ�7�=[�A�����,�L3�@.�`���,@Ћ��&������*K`I�z���;�2�'Z�Z]�����I34'����$��̜�K�n�2�D�n��.֗�ĀP��n�U�fM�Z�f���qv�]�WD:�����_d��e�J�D��R|�R4��=�-#���!���
������`�9��k��Ϧ��݁�E1X*�'�o-3j��C�o�e��;Q�<��w����v���m)r���6���_	����.y�L�ʤ�\͝ՇS��Op��(�e���9�k���r�2�Rf��l৾B5�D	ѩHI�i��Ж��R�GNW��؀`��A踝���_�/m
}�Ża/C!�Yu�����P��#�Ͳ�H��9CD"d�[Ƙ�I2���UeZ�@��&��qӺJ �U��Rį���:|��(UQ���.�gl��9rS�X�{m"�O���~d��*�Y��ai`c�h��'�L�p͘G�:֗��ve��6	T�3����&�L�GS>2EP�-�X*�B��2�߮N�7*2�T�����p��&.t�e�ؤ����?`���XKP� �ν��I�)c�W�Qa�Jñ"�IPqm߂
A_�,"�j�Ъw?��aY��>2/p�i����L������ÖsVM��%(v�0p�MS�\}� I�"��"���xY�䙧�����y���!�Mɗ	�g!�U�HGQ��=�$�/�~�]�I��ǚV���̴��� ��1���uC�W�V�<>c������v�;W�i�9��� ��^��t
�S)c��ZÃ6�ռ�]tvAT����$��J��3k���4����s���vE"/�m5ʗ�]]`[�Cʋ��?�8�'M̑=��s_��Q��_�=�N䭪���ڿ����+�P�dCp�L�������Fa���E��=�l=�i��|�$���X�W�)N��|V	Ɣ�T� ���]�[��Р�o�JM�J�׺j���3x\�W�`d��B�0:d"���Ҭ�X?_m��n�������V.B�5�{���aK�FJ;	�S�V�+� ��4�4�><�k4_Z.�h�������7�-�gw0��B�}ϧ���r1�c�I�Z���t
,[�*��A���J����B;J�--wd�^f�i6�d|���J.���g�]��G��N�s�⸛�5�����v,��<&���m��ď�PQ�E���3k�}!毲�!�* .0B�8�[9w����*t��Xo�H�g��`г�Wa��ş�C(b�����(�����Y@I�eR�MW[pX�wd/�9ErMxｗ��K�<Cu,��k'�k8�}��bB�� �d��V#\YjR |'�tS�5�������k'�����C�`dR  %ng _�l��}kBsCDTt���8���}�>k">�x �zO�ޭ
n+S���>�dɥ�5b��D��=�\"lZ�VX�q'i�k�yx�p{�>�B&�k�P���Ez</�:�a�V�ͫ���r�#dI+�w��e�����=D���w�V��Bd��^ւ��3hw|@�p�@,�[�*�d!��G��(��ډࠓ�/�{ҁR�����J9��h�0�X���q��V�׼�~�}Z'�E��G���Ղ�5+�W�.��#��;1���4	8�O���]�%C�F���a�{i_�g���ml��s�������Cp�,U7����Pb��i֮1؇���"��gw	ld�ՔD�������z�[N����Q/?���#�K��a��=T����+��Y!#����� 5�%����yF�d����uB�҄�n�)\�2���9qP'@V>���H?���0M�H��P@�^��#�7[������3�rܔūJ���v@�i��Ao�3�R5�g�d�1U5��
tLq�Di��'h��g�WR��,�2����V���W<�L�U_��bI_��i�oV���Ol��w4t/�ǫ�,��p<�5H'|�pI 7��\�1a�wn)���l�U-L!p�Ku'�)O������x���WmR�o/����M��EBH��Yd3ːE�1��U������V���.Ī.��B��D\ֶ���:��=����Y�~z.nE�4
DX���G�@s�d˽�	�fw�7����82L�Fi���x�}x�����X��İ�
�ܵc�.�nu�m���"؇5��[��^"�q���L�6�
���\C�����2`�>�r��#sD�N��\B��M��|ځi�&�{Z%HO��V�H�im��U��a�;=�VWl�h1�N��-�0������q��!ƽ����I��G�~
+\̽*yDbF<�=&N,�p$.N�xߐ<`LEC���2Z
'?C��o QYϢosr��~�+P���VB|5}Y�KoB+4��H�țFo]��r�Jͬ��&=i��`n���fŃ�:зN���/����Li��X{D��z_�q�'=�29�d�9x1M4����vE=��[�=1�9�Ud��\V�MN�{[�L�#��Љ?�J��!�
���yU�M:&�X�(�r֑q��iwd��"Y$yW�g�=Ջ���*E��ƾ���s	�P�/<�P��q����E_�L�#��T#� ����;�!�����\�u� 	JX�<$�]���grψ��RP�^jS��TK�P�'*��C��l�RQ��p��4������j�a&J�Ӵ�a{6�}����Dxh�9��+�Ȳ׮S:���#�M0�w�^�;:�K�b�B7�.|:<q�@z:ig<��_�t���S��87&�Re�@�D���� �cW�ǬV�E�����͏��T��3����s�+���[�h7Q�;Z�Yr��חy'뙼�}�#�+�q�Ds�Š�c�LH7������!;2�B%�5�� ��@~'�Eѻ����/�ۮ�i�j��a�@K�C����y��|o��O�U�K�qr\��eX���Ҧ�f��%|}2:�$�������U��tEr��P_���+�>56�䰎�.k���_gjO�2���,(�|V�F��`��+� K3�����Ъri���I���"���Z�mqӕςW	E�\?`U��?�ҮQ�>�0����xU�$��O�u�D�G���}�����6��Ωm�M���s�W.�)T����hC����yȤ/L���&�BZ!Ox�Img�^S��]��G+2[ىsmSO]f;�/��N�ϣ�%��h��tQ�C��(a���&%�>� r�ڍ�
���f>��5��q�v	�I�+C���e
V34���"��{����p}`�(ai��_����pI�j�~�����~�:�>d��
v�������k �˘�t�B���W���wHc'o�R�/z����Lf�ܚ3˪�j�{��ɩ �#����j���Gͭv]H�<���FU+f�v���]G�O��W��u�Q��?A^5��=t<��w�q�w��r�7�߸]�͘�&�1�˻|1���7��Z1���	��Jh\���BE>@��^���"A�1��B�Lq����gb���r� :�\����OU�%�jNs��&���C<���i�"�\�T���0�)�4���DQ�O㟐�@�����9ty34��̆���$q�6i��B���0u��m�S�^u�����p�S�0����B�V0J� p�:
�.0"���Uܱ�C���~�^����C��0�KV7��z�jX�qJ��������LyL)}�c��r;)fBJ��0���z��hR���I�4�?,⭂�2�>u
���3�8dȀuZ�Q!���< �O�v�sk%i��ύ�f��f�5
K`���km�:G���o��d���SE���q�Za��Ⱓ�[�/�Le���/�i�+�~ӳ6+k���9�}�
�y��/�߻:�Y��#AX�(#(4�A�C��@��'��~�j�D��O\eDZ��%�(T.���Ry}�S�~=2�����Q�N|� P�G�q��p<��������2}��n1�wNp�����ȉpd�}{��"./
�u�����lY�M�O�낫�/\^:��������PxR�x�������y��L�2�y�P�<|��&wy�K�y�pS,�C��h���vl��;���Ի��E�����nyVA��yp�h�]�$c�G���`�_T���c��imYNIl:&>?R��T�&�lR0�4�-@W�\���j%�)�>�͏��C�L�w�f���yͲ��B:qډ ��R1Lpq( �N�uO�0��w4����^�9f��Li����,��re�=��䩳3t��Hj�'�iD?rAu`p��"����p�!��-�49ׇ7����٫j��wC�4���R�4���mqSӦJa�9[�4��y��3��=�w,��6\�w���mrD�f�m&�T�gǈ���g��r/��3HQT�B ]��k�4�����y��67p�b�Ԥ��f<h�v���¯sM�_:��!3�RQ���5���5HZt��8V.��S���V�#e��.��F��˖a�3�>�<h�ϣ�YMv�ͯ9�hK�:�2�S�[V�=r��e�@��O	4����l��?V�4&�EW���}�m�.���U�
�դ���Uw9�*l���n�6�b�
�xW�3Yg���ҁ䪍���_�8��/�,ZIY�� n^�󶢆�U^�P󇑇�%��� �ޫ�8T��L�>iﴗr~���g�T�'��x�^�v��9uc&������$��Y�=J���/Z�v4y� #���&z�&�[�4�LJ.͚�	�'Ǚ ��<rԭ��R��*���^�HZ%Lg��K`E��������=?F��i	�5���oͬ-#1���$����ڪ���o�> �o+�Sч����+!�Ek�n�&נ�RS����Žc��� �p�����Cu��^���R%�H2���v�zȩMj�]ɦ�+�"u�5�_R�$��}���B�jw�H�f�O��0��0�q��A/�=������BA��6��#�$6�.{�t�O؎W�g��2�'�M��F�����D�ɸ���=S+뽟(�p}v�)n�7�\e�\7[+�o�{)�;N1��(�ˑ��S�l�6~�:��f�w��s!Ol8�v�o�]�����ۊ��m��V��k?#ۋ�'YB&�y�tGm�\�Hr��Lgq��!{��C�tF���^�(�e�⌤�(O��X��]�;��Jnf& ��!5a���\%�C��b�L��$"H�VEukOwa�b��J���/G�\D���N���,��*H����R˕h���Y����j�l-��-}��Z���8Jl+���I*c�$�0�g�d	zb����m1%*���c��^��&�lM���y�*/jDNp9�O ��``�H��FB>>��>҃ ��%
�R�]&Ԃ[#ӧ�w�dO��K�t\r\�
�Ǩ��3��$(��z��\�1� {��>��'Y�Y]�g�a/��id#�w~0-�eR�ћȌ
�h�� �^��K��
 K��k֢\�{��ĥߟ1n��������P"{ũ>}HP�����V/�|1d��VP���ׇ���C0���/��<�e��a���l9ǘv
�6��m���ߓw��[��]k�O����)J�1Z� .�SK��A\	��A/����w:���@�!
Ѩ�͂c�<T�P
��5Ij�?\���v��Fٜ?	�bPgd����Z��M7 ������Yǯ��*7	?���jm��񍜧����;�ȫ��g��gp����
6(J�=��
�;&��+�j�'���&���'E+&�O�>tz{�.��1��vU�snu�PzD+L����n���nొ�U�FW�Y���q$R�.���_�Kƾ���&ON����bX���C�u�C��Q�ö�3���o0"���$zk���,��y	K�����W�qla���� ���-��4���=���`2O��5��[*-Ԛ�us?�ە�k7�U�y����'Np��ku\�����u�'���C��O�B�7�~�2�#�?���������L�N�`�r���?�i�/�m��':���\%'qt�<�Vau��i��u��u�[l��l�+�Q��e��^�/���)��\N^���N�&\�R?Y�c��B9)�X���p�G����{M��S�۵(oU�)!�v�VN�]�n/(�Wx��2yсf���8D��� �
Dl&"���Cƿ�kl�z�fı���i�9+)����J%�鹵(�{���g�]l�2dI��y�'CA;����K��%Ϋ�f��!�&���"�Ԛ#�(M�����"u��i9:��B�۴��{5���&�IWKԭ����=D>���B���g[{�:QGZ�	��'�خ~#����4l	y��~����0MFy���Z]5K���6.���x��ώ��61o`[ޚ}���-].�@�aC�C��/ ܶxܡ
2��]p�|�;��v���C]�����`����G�i�&��Z����3���4���[�|��b�5Z�3-��k�:/��g!,��q?������'F>�xtK(�¾]i��t�"�@rJM����+��U���o�a��Pd��qdkR��Swe��7%S�m����k���<F�S�&�dH��&�K�u� �>���@*��0��-���i�xٔ3�I���v����L_.�hj�M%͐�i�`�M�� ��S�_1���ë@-H���v�a,�LE�����Ź#U;��!�p�0@H˞�R��'�Ye%��n0?>˥o�&�e����.�a�M��bB�����GKb�m=B3���d�S�`�[�8TD����͊��z�������x68z�Ӿ��ws]�JtN>g����+5C��	��V���#��TE7Զiz���3(����Cf�Z��VJ��t���B�k��^��3m����D��n���n��ߚ>��Y����@�����K#�fIV�}�J}(��	D_�����nh��l�f�p�R�Ӣ��㔍ع��u�&���zk� �BC���L�02���	"�	���C�W���4��j*ڥL��%� 5ѧB"!��EM�,����4VG����n��ڌ%-�cV�)���Sv�.^HV�CIS���Ð�f�㻓OBӓ�;/}�ɴ|<�������}����S#^?r����XБ��*�4�N-Y`�wD�jrX��w��W��w�V������m�Mt|����P��xA���
�&��PR�xJ�>P�ǵ��
�U&(�`Qtk4��An��v7Pӫ�}zo�Uh�qkB�(��C�aC�/�J��DjM�Hׅ�����3��ap|��9��(��x��KԻ��%e�[������)����E�����6�	��h�z��_6ߝXv���^3�#����Ӣ� ȓƉR�:�+C:Y4�;\�bk�PB<�;��A
�(��Vwe�z�n�)*\ ��ݦ»	��~/g�O��l�x��Oa��F�o������F��CS�8�ˋ��:(�3jM���*�7����Ш9��&R��B������H�/E8�i�˧d��2�)���8P�8�p�Z�Z>�}}���4B��������_��ޏUp�[�:G:�*�B�\�Kq
wm.�i��|�G6����q\Мá^����H�G��T�Ys�ݐE�`�
$���.�ޢ��	�D��yi���W|g�iɳ��=����r�S��ٵz��M*	s�ퟨ�����3���UJuo{�����y�!���%uɒ�(=/��j�ƃ�2��3�k1s6$\,��r�x:�S#��e�MR��oe�
�>��nZ�Y�A�j*2z������k��cO��{ ��yL�����=�L0�=��\+{Hh�YWbC���W��nJ�(���o��,��n2mA9-�S���P�w�Φ����	�o��ُ�l������6X�l�G�eڠ#t�r����Z�ǽP˪��ځoU�	��7Y����|���k�fї�A[�Wwyte�,Fb���WR�-���6��]�\ �$^:�&j}|xxc��"�$"�������~���䡩�5���eUǭmJ�*Δ�u!ҡx8�l�!���x��=]@U!d�2{��^Sv���
�;;��t1��ģ{�����r�����3��+�e����d�qH!3�x`�e5��[;���=���b��e�ܱ�1�L&o����jn� ��P_�Q���$7�T���]����u�cn�T3�ͮĽ���\�W�k��j;� �w�����|�b�K�8�b+�K56�Z�e{�����!�-���ʬ�ί��.�0�F��� W�A�^��%(4G�o7֭/��i��ӊ��G�Jy�Uu50�Tw���p�Z0�*��Mx	"�\��'M���j6d.�9�N ������Ti����l+C��Ǒ���zyO؛7��!��N�a��(ɶ}�v��6~�����?����TJs�0ކ�v�P��&Z�x�@7�Î�W=7�p�씯�2Fj!̯�b-����~��L9��'e�����7�?�*��G�=�q�t b_���p^��D9�7=��.�[c�Ϯt�-}<���}!�c �h�a�Ī�e?����������%��'' d_�~g͐X�`�Z�u"\y�WoS.�A_��m����ꩇ�{�CfbI���G��Z�3/� ��(K����G\��ׄU��0��InB[TW�(��=HjC��gL-�J��ŘW0F��:���,xVb{D1Ky�O���,C@6}�|�r�<����~�i(��p�Ɩ�4�y](2�k�f�����Uw�ME�r���@�F�!|��6Z>qY
�T�p馏ڋm��3�h��q{E�Tρ� &�����4_��m��,=3������Smd7�i/�=*����B�:C>�D���ߚ@0 ����-�eu!�w�#����eԣ��5�@��0籎6Y�:�,Υ�+�:~��{�7�V��B_e%���.��\������ٚM�T�:4��y��ϰ��@Z��Y�-[`�3�����F�$+4n��V� ��q�E�a�E_$wj�*�}l��ZU/K|p�RT�����DBveXHM)书����8�٘~��W��l��F��i��m?��W]*��Kz=�k/w�+����;H�+�6T�+�^�@�E��%�]�`�ؠ��
p��zϚ�kSA��-I��><�i9�f9���y��p<�D5.�!��X3����o� �*��-J�.�+*I���f�4<
�L���Mű�u'��Jyyh�/dreG��ڿ?nU��=a�C--���y�	j
UQ���2���y �u$$�dPh`5�Y�5ٚ�p�L���0��3t$U�Wm�����:nSqlo��eh���m���kr\m&[C��c|䯍�ҫ��o���_�*��8)��+������:�������_pô�P�\ha�O��a5n ���}�I�ɖ��p����w�Zt{}Qg��u��i��R�g���$aL�'�_Q�%�����Gxˏg���E5��m$Y����M�<���Bt�@�wuUo���y>��̠���?�� R���-���PԳ�N���p+����R��c�p���	&�_"im#��3h_虫иZC%�ݖ�j]bq*���?g�n�h0szܒ#:������'���%��	;��Ù`K\�<m
k����¡���K{�kue����y����2�1JT�sIz�����`�s���W����NT$���+�e1�ʂ�ߚ���j�J�K_�"��L��S���*��
%���A�BD����$�KEQ'�3dg2�l�e ށ��k�m����|��8w}H�����Hc�(q�`�ئ���t��Y��<�����O�m8�)T>���Q������IK>���ۖ-���P�M}��.�>g�[��%M
���z��8_���X9�Rz`"v\|ɐ\��u=ȯ�ē1��v��&|��z
�3��� &Ӓ��z�^�tpN8���Yu�F8b[.i�b{��bb�r��������Y�H媓k�pL�'��q�'}/襦+DTq1���E���[��V�
��#R��UwsS���=X����+��痰���޵Qh�4�D���T�f0&���f3��H�e�B�YfR�9ռx��x�W�Տ�
�X�B�;���»���D�@L�C٪�4���$:ƌ�Ø.!C��zgbp6I�EXӾM�.d{�aϓ$/U�(r������Dؿ�̃�c��1h��Dٮ��魸����d�aw���}���'��]�"!`�&����3n�:s��g$Gb��d�� �Nk^p	�j�5մf��Z~��v�Z��%���`��ߡG1��ǒ���$���o�A�xz<sv�M����r�@K����m� ���3zO�"�~{�կ4���{�L�W�:�~ ��Zc>W����E2�M��	3G���� �����Z�����R�q�*�G�
3.c|0)+�s����B���N&�~���x77oэ�m�<Z|O��ש�����~p�ؤ���%^�g݅��N))L۰�z��}����s^>��hgj�〚t�쯌iF�Ұ^e���>ŉX�������>P�s<���9��8��<wZR�#����a��!Q��Biv1��n�8��'��	wd���U�N�l;|���.Y�H%���ֿ�W�r?yM_�#V?G��d�y^OF[�_-� �V�6�׽o��Fv�Fy@���ڡ>B#D�6]]���������y�&�n	8�7�&���Ǳ�!���g�}qQ�l���QvȘ_���a^��p�6��&��
y~�B�8�V���o=(q"�7G�8I�O���a`ݝ�'�]�o`c}ѥ���{�L��fK� r�n� �rdy6gq�M�T|nΧ�a�Yäa��{nU	�i�I�'|=��wU�ۿ�o��0��V��-�沠ϩ7�v����$̩ӥwC���/D-��9
80�dL���_���(U%np�!bw��,o�ے�ٻ3.�����w���Lau-cP�i	[�oel# ����áUd	��twKr�=���1��L����pB��.����j-�u"Ub)���x? �2���7h9��b����Z��9ƲE��g��i~r؛�&=[r��t�j��~P.���G{�4�@���IN>1=�[N�$�G喂��5c�����H�y�2�}��2�r�[��r��(,'���H,m��/1m�?b���b�`0kq�4��>��SUI`����y��d���#��9��e��r *��j�׌U4����	8��%������B;�.R�ֺ�͢�dZ���k�E}�0��߱}�#��Q�6A?]�q�W�#BOf�g��T�؝a�$]�u3.:ͼ,p��K����_c�'�N�xM�����D)E50����
�f��!�c�`��r�h�.����#Jf��8CC�N�΍�I&s����W���^2�7��%���Ga)9�N����}'�8:Rp]�i���;��}Cy��w�Man��;w�QXEVn��}Jӗ���������V����ʿD�L��@p�����ɪQ9��4��t�V��RK�T+�.���a6��Oj���џ��q��[ lT�CA��D�����3���w����=�!7Z��x��K.}MY��
1���|�՜�����i��k9!ޕ���%�� m�6T�g
~96�a�ߟ>[��<��rH�'�v�ѵv�����	Nf�(�0�ǜ�I���	������`x%�c��whdI�.�Hc9^��I1�b�7�m��,ӜS�O�~7#���
��!.ƛ����e�߂V�A|�`[��>�t��(.D��	�:��ҐL���7]�mX�n"��Q�_��M�@�+ ���NJϨ.=&Dٕc��r��x�Ğ]�����v`�lf:
�'�^2>���ar:B�#h�2?��,�ߌ7��B�J(�'czx��La��ߐ
,��iZ�c��� UA<6� >q�ރ�;���ˇN�5���cU�f����߲ W<��������ϔV�]�όb�{�|�Un��������|�}ߙ��aQ�O#��:�����Y�YAUg��"������D�D��Q��*�B��z�2q�S5IﺓO5���=�q�!L,e��vy����ޏfgHnPi����^����'���4��.���SӅ����c�����ˌ��y���������W�ߝM�c�2N�p���ia��:�
��f�2Ϯ��_7����RƲ>t��yj�����6$:F}��~�C)�W�,��O'Il4����rW�쿜	"��/&l��Gic���K'j�xmo��-�*�SDyN�h�!cJA�����[�w@Vlt7[*�������1G�Xf��2�wÇ$�B��#���@}�b�O�ҁ! G�@�ޟE�؇�����?4��Z�ﮥ���x	�":�
2���/+T߬[)/�`o	�ێ�}�U
+LՎ	�=J����r9�U�>����`�$���\�ê����\,�û�C�˛DTO��u�	�f��8�&��3���v���L�} NH��3��l��}���%�qS>ua��ȉ��u$�YpA�W�u����b����N���o�4F��,թ�@}+�/�n�5A�Ҿ\T��,Du�{����@VЖ�}�u^ǯ��K�®�ZE����_/�p$�x�	�z����<-�"a�5�6���J�Y	};;���_1vv�����?�xշ[&�ܡUn�����p �rfUGEIh6��-��ܞ߅��2b��
}l�v���`�J)������\�5V�`�Z�#
D��/�1��	��1��-y��n}3�|o9�!e�Ca�v�1�/s #�Fb�:��N�F)��������l�SQ���D��k�� s����$�:�f��o�:�K�&m�$H�,�1�of�> �L�<��,�
! �:��K?�����2�s��MHq��	K��̑��uK��ߤ�j�cNg2E���X	@��$T�NZÐR(���`�sG�4E�8E_Mpz�g�TT��p;�o�4#Îx��g��@!��qIt�=��<���ӺI�ao�e,>�`�Nv�N���t�n�'��neN���~�d��r�B9��g�p��P|[d7k�*kG��7b�W�ə"��;�,�ޅR��8���0��M��M����4&���Ѩa{�"n'�V��������0��L����P�"w�����gK�:`�9���-[ �j[ *=�?���C�3L��2�G*Ž�w��Ns<��Gz�s�M��(K�H.lM�J����P�q}���⧓45�6�G"%��[�=�S+� 
yB���2�I�	�Qj�aIruӉ�ɗ;g��Nxҗ���֮��I�8��_��x���
Je��)-��u��V�6�D<���/9|�:^$z�e!�EG�g�� ���b�s�9���� ���(]h��dQ���Hyc��H4�����*40��u�,<�O��rS:-���܉!m��Yύ�k��S~�vi�k��u[+'݋=��N-��9��(�gj�jhým����O���D��bj_���T�G"m��O�䓑r4�"6�B����R�0F ��,��N�Mx�P�J����	uQJrs�U���$e�{�}L*}�d�:!�?Oض�'�X
��Y�i�(��No�c�<����^�����T�=��7G�J{��Ր�Н��/ĕ 
4@�׎�|��p��#�Q��Xx��c�����&�yXϴl������ݟ��b��S3|���3�k(�N7����-��!�-d[d*�h��c90"Tx�?~���6��Gd��"�����Z�m꟯oڲ��O)9�J�֥����J�X����4�Js�gN�EL�G����*K���a�Ev�^!� Q�V�#�yv��o�i$w�lg:>�B2Y������c*�f��B�+��ȝ>0�p��
x��>��	��rED����z%j(�J�?�$���F��i�Z�'�c���G^0���nH'	[�r�Q��+3��'��\��ڭ`QY�ր܏�<��6;I��m�ڣQ�p���Q��A�aqˤ��f i�jT�ͰD�/�|n��	L7IC��J����Ъ |��mD�✥ {汾���в!��ā\ �a	B~u�_��~v�H��Ɍ�Ѧ%�.�ua�\�q�&�4�t���q����G Xt�Y�+|��!�@N��2 9JP�!?i��b�w8��/a��_%)�J����r�#2s*��ǟm�����m��hu6�X���ײ<+*ju��z�A'����Ѫ9az�gM����Uq�nx�X��n��-�m�*F���U��4E�P`�Q�<�'����+S��	:	KI,P6(��p�o� tZgB[�f"/F<(n����2|�B�/<���g�sz��}R��*�H��F:fYd�!{����ur�H%*P*KJM���(��kȳw��1Gmޅ�kAܳ����<��J�Р��i�侣V�sH�X�K	c).�	3J"8�������q��YO�o��%����> ���5E�t�˳2�IV�mƉL����V���=6����$s	���M�WPE"����:U2�
tg�;�?#�gOI*c���[ ����]�1��6��
~9�ŉ	7a�a[���f=�e�K�hɰ�V���'�P�#+�.$�����[��9I�5�w~��Ho`2�nM++I�b�#����"ɑ�φC{�jC���D�ˎX_7P���/0�_΍��=��hR�:ӨgR�}!_�D��1����N׺��$�L|p���i�-�a7
˄��x��l�I%�d�f�4�����d�֩�ؐ����:�l�l8:�v5NIG�ĦZ˭(�[�č踳�\���c�aD���'��>.bQ���K�-����PY�2�.�J�3���r���闋��R%�Lz'�����"������&uFxE���>j�L|L��)�j�<~=�o�����CT�L (���Y`���wE�>��LT��(N��d��|J����D�.m承fo���T��=���y�&Ո��n��1/zVC4�_D��a�W+�1L�e�q�w���v%�=vWlk�~g	�ɾ$zW�∰�_�:(����2����:�R�9<��)X�cп<w)[�:%�7D ~��|f�*[�b!���_n]�)���&2͌b�����_�!�Xd�"���Fg�h���7������h�J7��y׾L���L����Xhv�N�D�,�H��1D2M#�z{�a
X9�)p�1��IG�m���=0s-�!� ��(���H�LLM�j�]O��X��HB����q��IV�t/�>&�Q�[d+Oe&�{3�U�E1,�#�BR>�! �� �3��X kp�&u互���f���;����֊���4�!���k�KC����a�֟�5��������%!�if(P��P�͵��N��rN�n���x4�J���k�HN�W7��ɪ�*�p>�E62{Β-7 pdL�j)����e�^ݲ:~����T���l�k-z�.��1:�+~_��wemcC�G�4���PQ�(YB�6yQ���_H�?��&�G�&�����y 8Zt���#����k�XR�C�۞��.��2�/�� j{��9Hz)B���Z�{}��4���0QÑ������u߽�&r�0���_w��a&*6�_���X�R+P8�wO��G�)������@_�_Q�#�Ji�&��{��U�j��Sȶ�����8��*>�G���?5il�B��Vϖ�Wf�*6�F@.�f�o�������ז�g羭����l�q������+��m <qJ�ZjD���{tzX�d��^����ۂ�ڐ�!E�2�2M�����C,f����>�>�w����I�2�T��y�^3��^��l���ά�
����l�J<Q2CP����T]ǡ�u��3E<z�Yҏ��}��.�Xe��j��1�üO^�zd��^������,���G$�E�hZ4��7|�h�>\������NPh9�w7jz�BD��W�l���j���0,u40\���Bl�]���Y�r!�E*Ù�݅�V���G��q�_x�A\_���`��)�&�i�W=hm��4M��k�r�D�� R˙�1�c�҃�3�wzbIv�ʛ���iaq:�5T?x�q���dpp�=���勻۾]�z��d3G�E�D�.)*���l��svj<~�DXz|�ؿo&�j�.P�xO��D�۾��Qd��O��Y�AME[��C&EZ�d��<!ʫ�Ad,;��Q�9�ݽf$�z�cnc�W?+莂k;`�4uy�?�	Yz7;��1K�/9�mO��8[F�^џ Y�=;qP�o�iqI}�D���)�b�l\�򏬪i^��jDd�d+c�O��F� �)����F��H�_}��d�r��g�Z��Ns�~��S�!N����7�xp�v����P`2_��O���S`��!�D��W�
z&� ��Ԗ+�/;��,���(qw-��؍({/e�����N�a:�M��F�b��F��G�`�����< �GM��!X�>��pI�H�?�<�S��֯�d��Up�{����c$$7��~��@�ZqM�R��O�	!���0������X���5�����+y�ɞ����Tx���GĠw����97/Cw�{&G&.��Z|�jT���7#��R���3��<li��_�&�?FD<"#�j�W�V�-���w;�^1-�GM����!��/��ؘ�ꕤvZ�C��޸�������~����p�nЈG�Rhi��`�[�2d#纞~��#�L���y�����V}��xx�(��V��~�"c�hZ�����QP���Kx��"9�z`�NEk��nՋl���kݲ�
�]�C����w�m����#�jx�>��3D�X q9�W`�XK�OZO�∟u&�V��}����/2H���0�W�	Sb�����-zs���6j%�7S2�N����9�$d��,���A:P�K��z={<
��|v����T,���'�-��!����p��}ɱh�C~�<+kih�G�
��Q�d��ƶ���Q���L%I=��	ᓲM������{A����1�(.�@Vj�Q�?���
���b%���^�q��)(5fq䁑�	G����d�+�`��^�������ޟ>*	Y:[�2�T�t�r	vc���(b;�pD\6H=�"����<egR��S���Өw���<[�z}T�F���\!H&ҳdI��ٕ;��\��3�+�q��$"����c�ҽ��G�B==��^�f:��Bk�+��C���ŌO��SSk���Ю���@>Ke\A!�oBِP�rx��.)�+�;吿 ڒ.�~D�ZB��0���W��
\����m��Ǩ�v�X���BH\W)2�2��ãԣ^M��8.-�l�[����s�V�尿���-?3l'�v��(��U��H@�GɂirC���zM����],9�+�K�P`�6�k@&~/�	����l�*k�N�v8��ȉ9��`$����;$^p��ȍ�l;4k��L�sR�@��Zs���?��W��% ��{����q���*�ڍ�P�K����nC��D1n�YFI�7��5r�I����O�U�5 yr�nd��,U[Nv�s3�z6E��Kـ1��A�3��h:!7 �wEz�&���5F2b�*y����8�
?Ô`���G��XB&4j����#������'���9_��G5/~��׏���RҜ���N��Wa����;0Q-D��;.*��}D�%h�Eϻ=w�<���pZ�ޖA���۠���-���U{�՝Z�dyi�K��t�������J�1l^ʻ�Z�S��~�86x��o %��-���`��e��aB�/� =�lKt)Gk�p~�s�\B(��&���8s���F��o��n���S�� 	��K��Lx��j�ϵ_��ʰ��3���k�9܍�|�ψ��&��^劫fj��|���b�j�� :��+{dcʁ� ���M6*e�5�'��[}]av��t�	r�F����6��l^�,�U�M,43�4�)�G(W�k�#a_��C���{Ob�ƍXz�/�PT�pT��=�2�1��q65jJ�ʎ5$c��,1��"��W�M��aP��(���4F�x�Y�P!���n{R����Y�Ax$[=�Q��<Q仢�,Ec�%?㎹%��*�"M*'��!0�/dH~%m�r2Φ!��ƨ��wv��}�6�x�~����R@�Z�j9��f�	eq �d	�u��^96��>���g�)&>�5|������� i�/�m�0w�'(�7V|S���i�y�h����>����d����S�+Κ�L�N}�#Y�+���ic ���.��2&ҖU������M`�%������^p"��K��3���������K���k)~SeuHQ%n/��gji�U��#���1����d�*�:�Xצ�P���O%��¾k�a�;���~z�
������?�	՟��R}�s������Ja���V��-\�-��~�wv0Js&����Z�D��໥��qB�S��������R��g�`�A^t�+��ԝͪ������-˅���RN8@߼��2�<��$C�0�?���⃬Pq,֤��:8^7><;h�L�bY���q��S�O3pj�މ��k�HA�y����2|�2Ŀ�������w;��}�&��K�5hB�㹟��>���s�/���h�oIDFPmO(��y��|�+������ G�Jl�M!v(ط@'�Ԕ�\v
e���B�m��^-���G���Ё�-]+���K#�q�70v<w?�U��8��������t#���<	�8�E�8mX�p��	KYh��S�I�I)~�Ad+g��ު�\0���(pS��QIl��
w#��R�Z@Xw�%M���M���P3��a��qlou��`��/2�|	����:�t�{�膂с�����}�t_��k��G`|(�Ki�佴��=m������,Ս��=�q� �g-��ܓ�-����G���M������{�S<������i�{���,$.;3A�TrM���&׾�� Er:0�����@�y�B3�}�h*U��%�F�e���0&Bʭ��oܷG�ҹ�B��*L
҂��7{m�h����?@Ht^�x7"��0��򚿀B�QF{�.�����Ӿ��H�m��z8F"�ȏ�$����Ub���[J��mM����^B]�b���4���!�$BL7�3B��7��د��ƀ\���z�|�>:k��g����b�/��ۀU;;�������w%ը�*�W�j'����Ӱ�DK�H�<�B�m����mv�DI����F�U�R�(.>��P��aW��|OHK�R�)�aM�&����$�P�Q��\-�������B/B���ܩ�6�ǥV8�>5i�98ZFpd:�Ӈ �5\A%����{-?�¡?]et���l�WO���r�e�L���a�dU�_LK�����0Y���?Tܸ�/�ue�#g��X�_����t�a�N�`KQ��������6"X�t�
����"y�m�C�UeT��0/�$�m]r5��W՞��L�2�V�4|y�1���0My�����  �3�#���w�#q<D��j�~�����4f�y�m����O�Pn�S�_m�>G$t�cճS'B?t���u�8�i0'�jC�[�L��R!�T�D�Fq�G��hc�[������Mu��I���n�9867*�b��±<�2c����.m�}�<�v��p�~���2�gb��H�#�d͡\	�%��]���AQhN
�����z�K�Kp�<˞�����$�6�V|�\�
�Io��\�3Y=�6H�;�L
)����S��Gv�PlU���+��*����P��0�L}@�� D������"��>�D�h�(�(Ȳ�<����R�Aja���eT��G�FT�D,|[�E�06^ �X�!T�G�Κ�E����Wؤ�7�j?�K������$��.�U�UQ��ۏ�kj_-�K>Ke�����	�"�Hb��R������t��)m�a��qr�)#�S�� #�r��g�O���?:����$$I���E�@b����F6�B6���^~�`B�fy�!�]Q�W^�M�ᡮ��A�͐(4B��L��$�s�x�֑c�������.L3F_
m�E�xw�EJ,_��|��V���kz 4hcZ����FT̞X�隈��:�ٱ��ڃcNNC��gO�9u����LW��Hn�������u�=�
�S�	n����*����ʐ�t��SV�.z��:uM1�6����C��գ�P��ǈMe��Ӆi���!y6�qS)sH옜�s��R
��&+��K�[��j5<S�r�w�Ф��& ��D��2}�Ğ�	
����D��x*"E M_$dX��C�R��&y�84jw��n�0r�G
�=�q+h�_��!���S=�@}�]��18���-�����y!T&ҀB��7	�({�Z�C474��)��I}D��o��k�='�o�u�4�Ǜv22W�8��0jy��\�N{����6�_�)�QY��r5�@�8�m�3�~� �)�s��F��ߦ���I%;{\�L( ,����KQ�_�x�Β��m��k/V�d;d�TN!�cy�vް=�si��}iC���& ��a�$5�ر6M���<pA�N��B�{��9����5�Svr��"�s&���a3g������s�3*���u��lP����c���!	�Aa�ȁ���&(��3�
I��WB���-�HҸy9����Ψv�����D
�؆�I�GaRwR'myp��J�T[��������̚������a�!N��ZC0+WN�,�N�;Z�jN$������`�Q2�/v�3�J��,k`�1�(���P�*beLN[�r��?�&�J�6o�u\�р�p��P��Q���:�0��p���S3��:��>KPV+[d`�0u�=���pa�R��L��_����AI�U�����"(w�Cj��6�G_zAfh�E�/e& +�'&�\���a@)�Ԁ��>�R!���;$���ju
y���4��cC!����,M�I#�����}��I��N�3���I��E�ř�c[
�t^wN$nF��SD�#���@T���X�=���dp�R+^��ܷj!�b_���1���j��&I�9'�I��l��DtP��� =R��PQh �-fR�"1�5��Tٺv��~�
V�zE�~�@�D�IY�㺬�
��a�ŉ�=�p'��̜�+0��\�)�KA�4����"�E^�!{�hHFA�e����f45^Hw<�֥���{%��a׈��������ͅ�DX/!]�K�o���|�3i����F����hJ�Tį�>��k�&,oz�6%�7Z�lΥT�J�C]��*�,�W4681,����? �*�Q�@fʷ�*��a�;�b�Wi����_��[���`��SS��]v5R���x��ݓ��բ��v��[ r���I�x��]%�� �ͻ!��0q�E�0�[�xᶜo�I.���?�En�f���G�5�05���y�tU�����dO���Gh�DO���3�;��. La��N��u	a���CP�J�$�ƅ��l���p<�v+�4����AsS&���)мS�CwLZ�P����*�]$e�' ѫd.�'!�����m���
򹍅�w�x�X�4�<w�\��j��OMA��(��?8ݙTJ�}�!ѱKx�2��5rc�G�]()����򗷑ܱv�KtY�Dl�1H��iV�����D0�pv9����|����`X���m|��k<.�(qH_��z$gF{�IU/р'	}+��S$�B�k��Q�l���F*�I��;C����"�����0��}h=�D텾ʂ���0���]�	����S�4�Z�O7�\�y^BD�"x�R��L�G<
�ZJuGt��H��H��ݗ�Vr� �H2+Gg�
�h<aÝ�s�ѳR�;�<e9��S݆ߊ�\2���T�m�(x���W����!Ҫ�O���Gc�{-p�p�u�'�'â�`4�됬<�q(�w����nA�dؓ���Ģ@Ƶ��\�����(���(��W�K%&��#����ƍPl6�H!��sG�r3κC�Da_��Wg+g��F�j#@Ϻ,��O� h�فv6fV/eO����1�����G���Ƚ,���Ә}�-�`20��w�G��%�VUxJ�@��`����	&]>x���>��~\8�@�f*Fc��h�`��U�z���>�Vns+�����t_�������A?`Bq7S��A	\��7LY�ɾ��C�bL`nD��~���f��2���?�g�:Y�RH^F���k��	��V�A�#z�ei��֞e/OD$f��ҋ�߄��&��!�^�"�Y��/"q�����LV�q,�+U~k�e-��g���i��u�>�ք�t"��Tt���̂CG���p;_������f���vƜ(j����X��3P�[x����d�zg9a��|��L8-96H\�65�ծ�r�\������t*�N�o^������[s���ts��l�����_P��A���p�S$?®f�K�T��Ū7������tƱ�ܐq�(U�-o�&�S����%��٪���W�F�k��߂�^�c�r��@v��h�-{ŭ����!��/YH/�R���Q�����w�վ�D��楠&�*3�Fs)�IG+Rj�3���0���(���"����{Vk��w���b��vVM��z\�E"�J���
�q��eS�L���"�s��g�t��2����#>y405un���5(��y�2@ᬔ�7`���$�����S�f9u��ae/}{8X�CM�]���Qn���P0��%w��aj���?�g/�c�0�d�M��qY^៉���7��\�AP�!����a�|吳g�n�G�s[L�h��d�]�a�Z%y�#5�-����W.|f�І�6�	A�k��%s������T2�A䞐7�:+ճ��k�ջO�mR�IE��=������f>.UP����1'�T�cb'T���p5kW�����z#G^��#k�<K��G��,!�o�n+��0��0�kwB� �vZ�\�vW�W%��R`@�A�}�]|��aZ�� �}�]?�{պ�.R~N�����o�;���a��:��T�3o�ȩ#p��]�B��n,�1���
�a� ؅�����܂�L�z#�KQ%��&�i��٦�֓pf�m���A��tb���jv�����"�=�1L�9�\����p�}���eBh����f�`<��2�qϨ�;�i!3G~����=!uf�~*4Ğ�<&x��EmT����*E��X∻3�������~�$����ﭖt��a,�s%���[1[t�;QC���*�ǩo�(/�Af�;9�7x�}����s3�Uq��|ϢB`���������$��
8a���0 �<x��Sǈ��>􍴭�E԰�	X!�8:A�	Vr��wk�����h��=t�B{ sw�h<��¥m8ۡe5��|1Q�I�od��|�BS�� C��Б��v��;������W��H%S0 U��*`c=�7�u%$5@7k0cW���6�i�b�?��Ö;��˵�w�����f7a\{���I���|İd9H��M�uc��dŢ�Aޟ_�AЧ�6d�I���:-�@��ތh�z��h8 ��1q���cscR����'�Z�9�w���`P�]�����W��n�F ~�6��|�J�?�	S�tP�j�fZl��hL����A�[V�Uxl�}��E��5U8w�2L�,B��`�u1��9Xa�{_��|M0s�:�;�~ND��u�����OT����K�$ =�P�»_T���]��62E�/�ɚ_�21J���!̰m�]Qѱ�@j B���,8��&:�d����I����#hO.Ӱ`�.�XPhm�	���F2��r|��/���Z�
����l������݂�^tB��8�޵�Sdf�|�n��;�ǷYA�P��|^�=�15�<*�w5�9"'!���v�Ma_-wP������h�dTֻ�"�c<>�- ���>��ũ 0;��2�����a$�Gl����x4��-�fV�)���	\����L��-"�i���y�p�e\�'T�:���W9*�k����i�����]u
���~S�ܑ�C�x�Z��i>ca�r]���8d��	�z��W��=, 8C>Oh���� ���O�[�.*�#^y.����D#�w,�����2Β��� �I�8�&����i��/ .�� 0���,�D����:H���:պ$;�'e�u�?>�������&�A�n�B�1�}"14S��7���h ᐶB�:���c���!Z���54(�f̥	�ܠS]��/i�P��A_sS����~��z�z� ��ɫ�˃�na,.W��e$f���y��# V�2������{�@S�8�Y�vgnATP&!i�SW����(;��.r�m,���>$ �i�
:�K�H˃!� ���NC��}�L�뮞[���cNvř��*q�2�JD��Zf;�~�.�)�`$�]��<1ī��S|��㩧�C�����a�oi�%l8c�V�pW��z�g~�%M�4,�/&����1:��%f��ƼfR�ŧ=t"�`0oR���V��3��� BV&\��1톊���G�׾���������
$wT�����n���y��ÏaQcY��_F��������[��G�Su1b)K�S�d�D��c�NJ�����r�6Z �B�Ѯ(U"US��TK�T/VG�Y�=�ڗ8:n��Ɏ�s���7��Zh�����4c��괪lSc����y�Ȕ��ϮԧȔyb\ʑ�<��+.�[�M0Y���:Y	
Ț;�o!���H�U��frV�T�ǳ��q��Wr���Ѝ@HH0��}]�����,��S��k�m\��:g��m�v�����ݘ��Ny*J'o���~��C�8�z� �%̧�<!�[0e�`�-2Cx�tT�ը
t���K<7��99�I�������>�k�;���1��,���ٰ��9�ݖ�pPftnkf���뒦�	a�`�h���[K�TY:+=�lO��Zջ��&�om���(��R�xi��`"U��w
(�z#��G2��n���8��4壧�H?�U2��ҐG�|E�2N�MU���>.��X�k�'��/�Pzg�AA�<0*J�Χb46�ᕜ8iC!��1��%���Lu���b��n�^��c���0um.����i|�(hϲ�����~�qPs%��maP�I?���vM��y�~@A*�|ϡ(�ɇ�z���Z�\fѪ��An���m�F4E�>��T8�ේP��11y�vm]�%o����Ma��#W�$��5X�m��*g@6'��m�B���9�/"��7�
4G������X����O�7�*@��%�]7�e�����M�:*�9=�r��
3L�B[�vk$!?�魚��2rH�*�[��E2�t��@![D�צ�������g<D�,k�=4�df�l�����a�!b<����]��?�j�����Î+XW(��d{:�swxJXb���ى@�#q������5u6E�ËJ�x4� ��E��ZӲ~6��Ѩ˗`>{~1���o@慹(��\ڢ�)j�`�qs"��9]z����lo����������'3��:�_#m�2����NO�?{ĐE���1�I�u�������G�>��u�u¤"��a���^�� POa�((PWfC�� ;d������bvޗ����#_���p�v4���[�TT{��QP��BhE��k-��X$p��\�V�򙱑<���ZTF��~NsQ�q23*�F�:�=M��=i�t.=L-mH#�c�>� �#pH�ʵ��{�P�J��R��A�V���gM�>�.�o�'謗�v="���xl�۫�tڢ'TP��Is
�x^��b�(��*O�g�B�;�(;��o��,BTj���