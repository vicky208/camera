��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V�B��&�8D�o��t��}��u�;T1{?�!��Sҏ�$�ۗ��&~�t�ji4N����頀w6��-W��*�`���.������T��ã�E�:}Y�&��T���v(�mL��P���A���Cؾ�n�e]X����c�08�� �v�*��n�s@
AgQIZ�#I�8o��
P��ɋ��|��e�WZ��+�%u;�$آ��h�xIE��tl�;4
�U�����sEv�F(��Z`O�{�rBd\�3�#��fu<�}��X�����BO�c���� lr��v�_��s�3�Z�����iP�t��� J�st���۫~��D�?����ׂ��>�;p8�L�C�&��ē�s�;�y�5�L���A_��^��	�t�] >5��[�<��0!o�������M2�]��
��ֱ)�H��=����<�E��^�^XY����y�a�c}�Ld`��e��k��-�؞�F13KSN1��f���n�ж�an3�3��n7@DB󠵎�F�	�j�y���'wI>{�L�Ȗ��(3m�D�p.E2�Ҙ�Yղ�o�N>�WIM�	+��i:6��3=9}��fO���T��[��� %�J�\��P�)Mc&"Ƒ�אE��+{ro3�
j�ĸL��o�әI��_k#�5�;���b�.ԷJ�Bu8�tI��O��S����-��$��V�5�/`a��WfaC'ው��V����/`CfU���}�
8F[Xȥ�: ���	=I�TBo>����G�a��{fQ��,������3��(ЇAɱ�y{�������p��;�L#6�fx��ۙ���0 �ڢ�N��$%@�����	Y\��/�6 �˅�������;��fQ5ȇ��r���ͼ�5�)wؕT�+s��\H�&,nɣ��[0T��-3j��pK�nL��Ad ������@�x7��߄]9�!�!���(��l��-b\�%��
���G��7ɒ�ފPZ����^w�����U�5kT�0E���  ���G둟ht�R����*�ץ�o�8�8=�� MGj�U�Tsxo\s�Sk�w\�l�Y�=+�@��ô e��i��|�tm���Ū�a��t'�^��-��[��W1�w��R��m����2�S�_�e�frD�.���\j��;g�6-t�k�<o�#�'E5��q�NK�����9��b��=��G��~��-��S��=ݨ�RJ���IKK��̸�s��7����ѧз���V0��V������_��6�+�5+�'�vФ��c��"�ulLN��T��%��j
�!��N�W��V1�� 2	6�ڥ_?9��HA��\���kPH�;YK�[5m��j�.m"!��l٭|ɦ���d�֓B��L���U W_�����l��HK
(�����U^/�H*�P�;�fRrs_	'�	?v\X��vtw����,�2bg�_�6��(�8/�N�r�p4D+�#���b�6����o_�y�������!=$�-�#*��塠��#�FF�.f��������"e?(�e���J ��-?;pс�6�J��A�Ĉ�r���Q�m��:���j�إk����U�@�OQ��S/fz�-����t��Qg�@��4��>�/��;+��=",s#����d��j[�x7j/��:'%�u��q_y1�ղ�H�R^V>�
~:΍۫+`$�TD� Ds�Bt��4��Q��Fi�BC�{$�ͽ�c�-g#�g��}�s�4T�Ҫc�T{�(��tO���T����8�˰B��E�\�s����,\�$��Xz� ����&ݱ�ok�E�le_p(�\#�[���,��on+i�1|S�8�z*����� ���Щŉ�N",u�ʶk�\��S_�h6�Ԑ̲(Y>�J�N����Z���=����Oړ0pV��}5�À?3*�.��b������S=e�c4�yz�����ϰ���0E��ע��/�+���hg�j	!���&�&��̄.���u$���бɧ��-�����
E��3��m� �L��!�1_��;�Yz�S�B=>�J� s�@�r�>&�#% <}�����yQ�Pd8��W{+�FU�2蠩N���bG*��ͤﲭ �4&�"m#�a��K��&��;��n!����;�h�+�P,���ә��$Wj[��_�d]�#`gb������'�Q�
ԙ �A���ǣ���Z$K��FJ��A�h�U��ŘK�+)��m%2	�C�~�!6����os9?�w�L�� /ᚩ�[��ť(�ہ�L�д;O����!gx�����ޯ��6�u�[���?Co���CX��1yX� �$����l�F\w����v�W �w�XuB���7�{J�v��ll���A���w�Osh��q���$lD:�j���d�a�],f�Z��Wh�%�mb�ޑ>qrѳ�!!�V�h���Gh��a>��=�2���/2.�I�,o�h�M�H��`hA��Sw ���1((���~�{S��=^����p�� ��_��bc	�aQ�z�u�N�d�SD�`oMtV.r_���n��U��#�����%�#�����0-}h�`�`�u��m?��a�"_%���j��sZ��ؓF�q������?�X�ӟ��ji<�9��YSٞ����PkqȘ�b%sO���(�ȉћYJ]���S�P�W�#qM+Q�N�{)m���'��L�VT���W�oR�K��
A:?k�zz%!�$��L�����S}ڼ��){��̴����*�@3r��SY�L�Rf���qR57�lXJG�B����?��*�X�4���'���,�rD��7�����<��K4��l.����".Z�'p�qKp¢�|�F����|����@IE�?7��3;��T||\�b}Q���M�U�^x��#�~��f;�-�|?b��_�	C�'ˠ���{�o��rߥF�Sp��V[���OW�_hi<�M��A��Y8��n:7Ⲻ�YJ;V'�t��ڋ(,2��y���h#��jn�!���[�f�#���뉾��W�	YY��{NJp�R39f�,��*��k繰�#��%)�5�!��5��
=L�x嗞C�^6�L�����?�Յ�"2bZ�>(���w���8&�j?#R׍����rD[x�(�Wd7��9�y6�ᤊ���2��f�DhO�n�q���c������ܶw��'�ț��t	��w3�gv0��L/0@+;d;ܩ�Mq��;Nl�n�u;�iJA�%��?�f�>b���,��D�xǡs�T2T�j�;����+�X��A��a����D��=�ĤNIRjW�h���D-����[B<�f~օ��� :
�ꡌ�0cX;nt�		�V\Xa�k����K�c��]�*q�>�Z�2@֖�K�ɶV.��w����)q�琺߆޹`��0��g�P�͠4�Rak���lYsv�.i��gR_�A}�p԰�D���V]7h5�U���tn>�_w9P��ʹ{�����'0p"�R��U�8��?^��a��~��%��3#aR��[`)��o��Ս�$��6���#���UN�8���]1�C�y%ٓvN�\a0��X��*��
�⺑ 6�ϔ������m�Ê�à����r��"��=�3F~.n5����W2i��N�����H�6v�����>�Ϋzz|�x�%��o�.Ym�O�y�)����Y�H�cg���g��q�$"�D������2�g$���o�H��6�-�n�<����ALk�}r����q�3Z=�L.s��x'��G�q��?>����Jh���7�ܒy��[`H&W���V�Bݰ|Z>z���|9*�\U	��m&V}��}���lS�7ʼl�|}j?�I���^۴2 u�è�B8]�j9�����*���	u�=��оR�l��[o{�9��q��XF�n�-eEp/��U�т���`��$щS"o�78���ҍ�7���46�.c@=���o[���sQ�	���tW�E�K̍�m\6&�>=����j�䓫��$�~L�	��*<>Xg̠)%��|"_�ܳ�/��{Bq���[�9���/)��|�,lz#j�N�&m�S�ШhV�=\D�q�PʷQF�{���̀^G�  u�hA|#�u��Ti�¢��`�m�e
I�#�T�A�T���9���G�XhC˳F/�<���i3���RB*(9�����}��\=wB/��M��[�kȝ�Y'̙f�hB9v0��g��{�j�|({hOkT���OO��>:�Y �1�*��P�����C�v�j�~�E�a^H�8�,LC�0�$X��r��^�J'��\�v���Ȉ�|Fh?z������X�Q(6�#������+@�3 ɞ�4~�0G�:�c�Zڊ�ykēU,1����׳�+��\նa����W\į "¡���A�0����Bår����@���N��)Uk�am�6�ck��_��������3(���A��:�CѮ8ؑn�"�� >��uv�%�¡�E��Ŭ4���ׇH�j�a�&����d�!�����K.1�E����'.�$�l/6☤H7�E>��$�ټ�o��؃��[����p��:�o�C�՘���9�c����+���'��w����ge5{b��(��$�R򅚪�1���o҅~�2(	~���~O_�]��Y%�sJ�|q9F<���<)V�&�;��w����x/=�����bM����,������o�%��$�&;i��}̌$�E�0O��{7��Y�2������(�w���|Q�*�(%f�S�	ȗ��`�Lm���MB ���K㓎���[�A�{b-uf�p�+e�)���|،,G�Z$�ړ�P8��ٖ����95�?{���Q7��(��"�
LOV�h\#�KЛء�1���1���,[���n?QJzE&�D}�u]���}�Ï�|�(\��I8��ִ$��q��4>��[۪����?�w'�Y���@=�5N��ӻs�ٕ�?�P��r�;�az������b������>�K�[@V��|z�N{�'���ÝyZrJ��h��	f�4�<O�0��A	#`��w�Q���m�6�nĕ��,����^H��C{r/Ｖѳ�뀕,F�m�>�Ԅ�sc�{�G�<�H���6��[�����U��C��޳�4��XA���TJ~��N�C��/@E}�-�͜�S�c?�B���[j�=�]��(w��Ա�*�LЧa�"�WuP5ʸ�$��L"b}�sDhS�uF��.D�R�N]~<b���h/3��G�޾a$`1�.���W䎉���X�pT��RM?1�g��t��_�ȵca��#R����|A`������OD�w8�]�2��`�z�ո�Jы���C|�}���}��w�jg��r��|�7L�"�~�߿!8����Q��A>&<M�M���Hn��V[ZТ@��1������J�_�������ָ��۵Q]H&$	�SZW#ţ��Fc ���K1�xi�2Y���S�Ng=���Kݩ�"�9�$Vu��M8��Lؤ����}<��u��coQT���A��:�O��a_Eʣ.)�u�^���]��F��Y�JEI��^N&}�� �K>Wv X��� �����(��aJQ�����@��ɘo��"�/2 ��zeVՊx �|[V�X�3�z��a1��?�CP���+���,R� ΋_����ƨ��_ݮMǖ���uU����1����"6pw����|n�/�7��?Uwh�a_*��?�%I�p��Ez���y+҅���4��]���}����O�o�g�8zX˅��S���F�쥈�[:�o�f���rm��h�ĝ�/z���EV���:s֔`� F���?�-�/�`A=ES�1֙���i�D�*��BU";X)Y~f��
|u,�m�I=�߂	;I��	����(�-3�Z���c+j;�_�Z�n���]�����l-�I��(G�c�08`��:�z�X=8�������.���3$���wg���L�l�|��Ɓ�/�w�����4_�MZ��a*�.�>�L�;*97�H��E��:`ư�%�I�d}���n�w�(C�giG���)�顽V�;�+/�E�8��8�O-��T:kv�㟢�S�YG& kc8��LɄB���>��1Sza��?�(��|�*�
��<����6(���*j�������y�	@��(�\npinhaA�BY�~&DS�a�1�C۾��Z�HݽiU��-�7���>��O��[5M\Z�$�O��FmZۦ�8�k���H�#C�~���[�S�GpԖdp�cN�I��c��]cuJ/4&���F�U�x��'>�r��0����`>�;��>HMZV1_X"o]i4�@Pz6���&�1h2#�5E����� � ��-5����)��t��2�^�}<�4}�ݘT)����P�^��QJ�~N3�i3"�^��ԩ�; 䞆v(�Nѕ_c�]��(ch��N��H��ƾ[��&݊��q.,���3M�a�80)�v�>n!�87�Z�@�Ө�9��s��MY���������o�A)х�@���$<��;?LU�{�5��T���D��� ��~��\W�7���d��;�w�e���>���3h/�U��C�T.�����6���f�`�=wD�/Ν��8�"s���@��Aљ��(vK,\�b�jNئ.X��7R�7����ie����Z����-���Ht-�Δ[;��<񅀃�}��$\��?�x��)jD���Z��],(�0x1�A���mx�X�
zm�m����m�_V��{'�����.�bΙ����`��U����8p^�w�.h���}dy�����	�|eq@aM���bEhOKr�qԸ
4\�Fp�|�j��s7�Hܛ@[������m��8�R8^�k����
e�6�V?�bK\��V�ۃ�w�k����4�9:�ŧ`ө��U�8��ˑ�]R���`ݚu���Υ+:�&#�G̯����g����d}�><M�q�nR�5�Z븃�M����	���-�U��]>�{���>,O=��;[�0~��T%�
�C�R��:e��ѡ�*�b�4���ӆ���$�T��:	���ɃpD뗡,�@��d�G�������M����R��(Rd�z�ˇqy�� ��ukkTS�q���{-r���y�^@�/"b{T�ӱ�^1���Jvx&�ϡ�.�/�Z6�W˙b�_��Nv� t��H�Z
���.����^۴^a���������gؙ�G[��u��r�p݁o�O�[�غ�g%�C����_n�L�_�b��F Љ�mw�RK8���<�)�$�ٻ�b�E}��.�URCW:3�dG<[J.��:��2���{�]�hd�k ���N��2��D��i%H�v�f�:i���NXZՇK$��-�}�����렅��,�٪�\B��:��#��zC��
i@@��Tf�P>�V���H��ģ�=_�v���q�����Tr��]T�K��e�jF,�uFh���*��47��?1<��ڐ��i�' ���JGFE\�������tu�=�X؇G�8���P@�X����:f�0or�d��y������ÚZ�#8R��ľW�f~��W#=�kw�.�3ǻHz�6�~t$;��(�̲.��i�Z��!D"���pN!_�;��H�C����l�ػ�d:LI����ki�Q]�z��t/�vKM	Ϗ��[XS4# �Aչ|ޭ��IN��԰�t-$:]N 4�P����{/ l	x�F;
mK=Ck���c�t?��\�f���*�D+K
�cbj��
�kܗ����E@�b�-d?��=�>���:�j̝�If?r��P���[��.��3�+�	�7�-�*R �9�L]FKF�@��~�yRÑ��ܢ��A�l��hl.���x����[�*�ˉhO ����V^�d3�^���o[V��|�D� ���@�ky�aZ��\^U��;ǔ�	������-S!2����K�B��4���g�����U����rgG_Dw�k*?$�Gz]��+��4���ćw�l��J�C�(FQ="�W�P ��~�@>Kl	?�bM�`~�Rxek�v����#��V����Ø]
=8��}@H��
]<0<��!������l-�R�W/9-�Po���ye2/߬���n�0ޚ�}<	�
����������Rt�5��{b�J�*�!�K���^�~q��c oZU��w"�!�sl�?�I���k ���F%s�Z�Ͳr���zNI�Z<B��,�5�����--[��W�m��j���X�K^�#7�&�S�߃qį����?1��da�Z�b��-�2��m�M3�o?�d�"ʪSP�:�[�,�E�A��B�Uu��>�)�bq��7�S ��!b׾���vh4�x)�b8�@"e�@f����Q�>Iq���^�Ԅ�c��m�օ�>Q�W��M�(��kM������Afe���'ج]w�P���O=hXY6 >�@r�rF�پǔu�B����WP���8zfHq���a��I Z�E~6�E�}%[Otv*�)N�TN��*~ 24�5痧'8xr���+W�!�c��\2�繌�����.(�⋢q�%GH?@_�\�ٖ����B��3�;��ۤ��U��qM���-�e�<�8�������ԁ'�UH��\�J�d�,t�LfS��b$���%he�My�1.�F�Ԓx�b��QTC���3X:�mNt�[[�M���\�ٓ(�1J$��i�Y�M��;��Q��Vo�>1���ñN��&ZE��'�:��%�K7�}���)����������9y#�1 k�q��%��*���)\M%),W���87Ѫ/T�c$�w��ϯ��@;�sj���6� ���Twn
����.�"B��~ש�;� ��q0ۡ��[^.�
�C�c5�ê��^Ӹ�k���8���a�խa�r���;�p��d��Y<�J���ґ���5��T"�Ъ�W��N0$�K]4�T%�v�U��չ���fІRw�=XKM_�u��#(���2$�	Y�v|+���K��
�����[5��c)?�d����:^�/1`O������7��Dv2�g���<q���ZN� �R(��nL�Q�@g:@�~F��-~6���-a-s^��\5T}4p��$X>'�H���ɥJ�c�fu�7(օKe���ٖ4�N����YVT��E �?�TNO^�ҷ�G���p7s�'�l�)�;F�cb/&qh9�'=q�cv\ �4n���+�8��`�T''teA�,o�8�Y�@
�k3��b�ʷ�_7�g�m��\���C��,�d��s�NtE���Ӱl�d�#�e;�x�%Hۭ�s����پ1D�G,�2�:Ɂ�ƽt6i�����8G�����.� i@8��!���6'�k⽅����m��7w_/2 �;U�a6�:<Օ����#`���Ͱ����o[Ԓ��`a�v�y�n�;B�9�>����ӼPw��A�&n��5�a��fu�ƕ�dg�u'�Ŵ�U�׭�d\��\3+��e'�$v[D�����d9(WT�������C���_����*������Z�N����ٴB���8x���]W�0V�vy�?O9����`�;�ءѼ�N�]ԯdGr�����I�>��ׅo)z��yЮ[����~�����v1<1(�C�ũv!��G��<o�@��:�JfG�u���:p��(y)��i>O;ԋ +����?��ȏ���lCE��.�����v�i�cA��E��4�,�)�f�a�,��Sz�M�V�筝��	R���X����Ec��>����H=�m���:j=��m�3���f�6'^�y��u�w3|k�F�B�d�%��ߐ�j�l���fgOP�'�]l���v�q��{�|U5�g4;E־cP�`A��^�[�'َb�r�������}uT�����=\�8F�oa��YT ᦙ���6~�n�]����2o���JC</@C��N=!�������UW�/�_�hQYl6�c� ʉY��a~�y��TT�~Ï���Y����5F�H,�*��M(�A�4#,y9������h:�l� ]^�N��r�dF���Q\!c�8s�ֹ5	���=s��V�Fq�2]UN7��*kN�K(1�A��dW�����2~n&�R(�(-W	�J��H�|�!��:?���831Z����3E��o��ӓ����&}m��b\2�E����=�r��j�5��4��ax�@I�m�˂-����\�ਕ���V2~)�A�<�>�� N3T�`�}�~/-��[��|���[؛���.3��|�s釪�'+�"����-GN�Z��OX���^�}�C��+]��ql9���h'Ւ�Tk[. �*�����i�%���N�I_=�
b��{��r]^�;X�M��j�A�� (xTS��i�(�����d)S�\n	}/�Pt�&����#�ypV��+�&��ԗ�{��l�$V2�J/u�n�7*N�&	��ި�D�E]��"|��|ۣ�:�։C��>��,��w��-+���A����m�vF�V}W雩UP܃��"d�{xEK)8��FT4ʫƸؖ�p~[�-ЬPO�(�\�3���k�3n-���L�뛩x' l'8(k�@./=��8 �b�B�	M ��I/�9M��[ ��Pź+�?]ٗ>�����]0��h�?���74�����<�l�RI�!�aT�^���&]_����2�� -��X�p'�)�̓5�Z����̍��������~��՗���*{��<B�� U��������#Z���#�W�����8����,ϕ@�&3��o2?��gg �|��Tk��M�*���jKGD���hH�����p�2�Z��Q�w����^�Kh�ѣJ!����]�`Xƪc?�z�0]�@@��)Ro|�g�d��V�\�ʶ��}������1D�.�b4hAyG!��	W��|`$�@1���e��U��<��W�5�)��5��b�R�1>rOhb@�>{'�c������}�Z߀��r���Q� ���S�(%Ju��q��@���H��>@Q���~�f�z���^��.Ź����I�q�颃�+҇��V�a.�.?Bʡ�7~l�H��^��t?���>4������=�6�v��_�i!��!�0���|o�ؗ��a�5�U�M�E,�I&��`��t�R����";"��j;)�Q3��s��%��i̊F/vX[�$P�i-$�AV�F�/���[�=���3Ѭܵ�i�Ō?�	��{]���N��[;���ķb)��.0�9c�Xr��y�K[�ѧ������8����S	ˆ��G�uEO�a7p���FI�=`����R`9r�xt�� �_,axK��MZ���[8��{���`�G<{����V��A����>����V�V����<�n�Ы�4G�rR:�yS{�#d�~~f2.m��px��B�7�[�gӤ�d��h����!�q:��ɘ����f6BmS<ӕ�����݊;��b���۬�C��2:����E�`�)�5؎�f׵���3/������>!{����_f�E��[eag���Ȯ�I�7�X����""��iR�� D�e�+?��򠍥@&�K�&�'���U�6Dz��d�3�b�ߠ���Ӝ�ķ1�ZIV?uń��i� �&����jg�T��T%�Y�*K��l	�)�*R|��s�#l+�9�K]dD�W_B�+����z�.���z;
{�+le�+/�z<�h��.c�H�ɳ�Hu
d���ٚeZ��H��7s��v�}6�5����}�Ę��q�� G�ѼU���h�n�eQ^;Ov��|�b�}`Mz�b�쌩#�#o[���.]2G;���SVQ!��xO�m��?S�iܐ�&s$a����(�FC�|J��A)�\��¢���Cy�\E3��Dm�U|*=�y�g��t����}-�*�U�*,gɢI�`�va]���d]�U7/ z~3�G��)��:�P�c�z���]��P��H�(�F�	n��^�FX9��;C�0@�QGr����5X͞�	-������zfEL���OJ�J�}fU��.7������?���4��ƛ��S���x=��G���������B��N�x�R�C 7�L��`��0��t�B�T�Z�4�
����(|���=��0C�u'+����ӹ$� [R&x0e� �(!E���$���4G��J*8���s�Ʉ+�Y��i���5kEe�@x�Ӵׇ,��6�=����M�<8v�hOo�Z��6$�����5}�ڥEf|[��5��CQ�ZP��ȶ}�������%��;-�A	O|]�����N�@d�%=/j7U#���d�aS��B/��AhbY
Ǐ�X<Y1�(zۚ{H��X���i=�;{j�*Aִ7<�F˫�Ji2sFL!�U���-��s(���o��3�+�[B>!e��aZ�}(�	�Ċ3�ꚅЖ挬K�3�#��*�+\�iΔl��8�#Ol@�n�
�7h�16\q�I��5g�d섖��f۠��J�I��fkXh�@�32�ص�2���Yʕ�5=�T_�]�q�� pVK7G���L����8���Ŀ��D��p^|f�Vr5���LM�	���f�Ԅ���_�Q���/�78����ec��s���-�h���~�jޅ�^Bb��L��p������Ʌ�X\�+�i�b��	�Fm|f�g����(�"=���-�M� ߗ��/ｯ�	�*��x��Ts��넪�{��0|���I�s?�+�a*o�W�L��G\�ξ�m�xh��-����rG���h�eM�$�-e=���r#��w���,�$�Ȃ��?#bQVG�:ܭ|Y������+���C�f~�6p��PP���a�O�|�e�����Zzf����م���f�UX�H��^K.{/�\?�S�d�+�k>������;��p_�[�)B��k�?�7X��
o��������Yv��t���hʦפ_�p���J��G��
�͚ܒ@0�HW�~<v�1ͭ�}�o�Ң9������$5�M�g���C�Ig�qT�C;�OX�.7�n$�9T샖ZǬ>&rB78��
����颿]N� ��H��m�k�8�up;5?}�T�v��9���ɑw0�'F�_`�P*}���
�?u`�S�3�W�'@ M�ҷ(4�Ă�q��Y�@��QX���ה�^��G9M�NT���g����O�,��/�B�'��3Dޘ�6C�?T$�T;��I�|B�[����w��<=�� ^�N���M&q�[�!éq1�Ʒn�6���QG�;f����56�)N��s'�N���k��pנO��uDe�0��
e�N���!8�k�v��I�eC"8r@��E��/�$�M6�Mv�y�͢�o���,dO$>Z��+�6b��<�� �j�6M�=�*<=�P��eBRI[L{]��Aj��Q"H	}��%2rs��99�B5�\�X��*�D�/Î��̩+ �Z��I p����?��@o���������:��q�o���sd�7��X������"��9.U�%6'� ��!}Y�����b$x(����UED�*D��E�����E{��DdG�<.�S_�sgM�s+�P۲�F8�t7�%*CW�K@����K���Һ�0HvO��шKei��7���*}����p�ze�x�h<3��gܝ���+`{�m��*�iq��7�U����t�� �~׿�Q�� �Y���O'�!�:��8VyQ�j��e3K4��N�lPeuDʁ��p�S�l~-;lL��~���$+�����q�/
�U�t�z��(�J������ۜ��%k��p@���W�9x��[���c9=�0R��F%��@z�c��L:��m�p �WA�5�--	�tI��[╫����=�>����d����u��XFA��U�|���
ͣ`����;��Ot� Z�v�: Ed��/��ߨ�K���C�/V�u��_�o4������֊j�v���l�t��#BST�������0�I|���6���1�����0{�47c6����MΓ���M@8��ҧA�)�}:�x���ϓ"�i�� �<�*H�}	�\����!Y�,��1�0��^�m&�YF�!X˹ʢ}��9��A޼k�����s�9�z�:Q��[`�Eb�RϬ6�8�r�C!�
tbxTJ	��$�]&9:˿�63T;��d#�¹��+�+���L�x�
� ��4*���C���I{y��&��r�r/���V�3���ԯ��Q�V~�*� 2�e���O�P:�_��n�N!I���$*I&�Ms:�l��z��͇{I� ��E>Z:BS04��� j��+!>n�8t�>�S�Bbr:�����������;����َ,�9��r�i�\&}�&��ɉ�F�7������0��!Ej��mH�\�G��n�5բ�3��#	�%J��T�Ő��ߤ�h3ӗf���(����.u�s!�����\�x,�|鸖�@��}b&��H9�Ǎ�/��tJ���	C�S���Ne�`�^�B�{���.�y�������7��t�I��!-a=�i�Djlh�[�.��8�����@X �L�<{0�:-��?��qBC��'C�uߴ�U�f�z+�h
N���b�Q1)����0���k���:�g� d���<��
#��*Z!���F1�$0�q$�@���C�[X,<����0X�kV��<�����m �����7t���_h+B���6X���J5c�r*p���74�k�nW������e*}0d�,�v
�D*��3T�k����<8|e�C�;����:�(-no�/O�,�*>�HP���*��a#�D�}TM�:?^�b�r)�v�e%w�9$��SZ;-��Zo�������(4���_	w��7��P���T��RDȉ��#4��[��TP$�yZ��M�O^�@�����.��Dߚ����]>TaO�ک�3�o�_Ly�ױ���2ś�q7S�	���#٣�³�:3�ȟ���j-r�ω�#A�N�
����`"��P��σ#�y���nZx�� 8~*��_��Z��c ��XG��ˋ��ˤ��Nv���ͱ��IC	f b^��`#�f(��[C{�	M�ɐ0�P^:G�@H��a��m���,S�2?Z��k�~݌DN�2�.�2m+��ڣ=�z�w��k���eb����k����{R��"�&(8�u��4�R����N����K��!b^�RL�hD�"w?,_TkLݢX���Ì)����i�"�p��=�9宾�z�J�)v�=p��G�1ᆔ�,�!��79�m�[�$�݅/��?KN���m��[z�*/%�a��.f�{�=3�\��%#��zO��M���DAY5��!�{�5pZ$�B���3�����!��)yʘ� ����Н�zL�C7�i��lb4���$�6��f����Qy?�� N�o�hXL�j��O�l�é��>���ꖕ������;�UD#X���\ݛ%T�i���$�0�� � ��o���Ea�+x{{�0��0�(�>0}�A�P: W�Eˎ�)G=�V�_�E�"��|�O�S�%S"`���!�bj������v1	�S2@�Z�40t�`z\���bp}S6݁Aw29,�
�ѫ�T�|���!�*�rD�v��$�|E��@�O̶1]�1�	��U�����b*8?��g$�43�� <�S��R`E��]��x&A(�����y!��G����_��iOw���#�<"Bz{�Z�W�7�}�)�ւ�庱,P�g%^h@˃�Pt�J� �4�*���2��U n�Q�j�!�(��*�Q�l��!s��qZ�3af���=:���#��KGi-=��~�}N%y#ĭM�O� w�}2��7�<�J?����wi�W��`��8�|�m���a~���(Ox��X4�
}��D���L�bʲ���;��5.�kMr��a����bF�c�nR*�j�c�X�!��9j$sbs,Y\t[S�-�=�~)�T���p�K�c���s�j��S�#�j�&���DQ��}S���WS��.K�qZR��AB�j�r�s�Z�kX�-�QF�g[b�&���~	��[i֊�t���Hs���u�D���=:6
�T��y����2�(K�[�s[0�z�!�i��)��L��L�Vi�0�[��.�,@Y�� <����f����5���CY��\}Iu�F;�6��9 K8�DύM}��Y����k�-O�O��