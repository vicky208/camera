��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:��r	���cW?5���%W�$X3��΁��P�@&T�V���a�����W���afDi h�c�L��Ez㾤|��������*���D��B`���/��8�Ѯ�'��1IP�i�fp���l��:��?���R5J[!�]�瓥�K��~�3�I~#������\�]p1_2���$l�&���:�ly�e�X�+Tv���T [��Q;����H�2�`��F�m|&r��|$l�ao�̖r�!�N.L��BL�`_�˲#�Ў6�a���dl������
|Cl�pn�(���������/?w�zvVH��r�Y��qN^r�'�qI|�T\P���6��T��?i���E��w�F����2��f�̝��BZ�����!��j�3���+��a��Tȫ�?*N��#c�
[D0��╘�쟷w�0C�A��ƅ�,�B�-t�Wӫ���V*_��N� ��<	U���l��+��������A���[�G7����j����P?�|�XJ���<O�r�X�̆��2Ǆp��q:��j4/��戡s�v���m*�^����tPh����e���}_���SYzC�x�zlN���l�k����SS�C�%�?g^ӽ����+��	g�P�V�"ص��!�:v/憉����Gar�r�	��Z�I5z�C(M�+6�{�K��8b�([:cR��Ar�t��=�=ݻ*�7���y��x��~p�'�OVQ��"\��iD,���@�����~�1���
Dҝ��|)p�|Nߘ��e�{h)J�/�\�DOֽ���}5+~�Oqݦ:�0�)�EPR�j�%)������1��,�O���5���|�l.�6@�rslt ��f�X}�~"jn2�W������"|��:T�)_H��,(J�6D�;zܑ�����������I�� �l{������䇷'$��̼ƌ���@.���n�z��"��4��`3@��d�=����o�c��{���@��@ �b��9�q�5����Qú#�=��jxKB�G��nL�ݪ� '�=�/
�����7��f�eG�`[s���C@��xހl��n�h(�}9�.��g��K�Gu�-N_�Q0Hn�Z��,d�9��yL�MR�ک���-
���y �Z�		g�����=�^���ӑ�.�
�N�i-v�y#/�n�@^�w�%x��V;�J�3pwC1�(G�@�'e!S=�B�q�|9>#�g�Z��_������(�.�lU�f �N�-�;P ��M��a�j�&�����^�y]0ޠ����k:��$��$���w���u!���0.#_�]��řB��d߿Or�D[�W�`=���Lq��o��_w �$��׋�R9�x��{��MJ��ٓQdv�-˞���}n����b�I�)|a�
����HH�kA���VU�G[<8���ǩ�EX��9��8����g7�ЎE��ߘ�/1���v6<�Y�J�|Cf�=P����*�����ͩ�y��γ�/�s)��>�7�_�.�/�M
�& �&���7��:m�14�v��'%I)J9�/<�� �B�p�n]n�J+o�,���0{`4a��P����§3C�Ye��I9���~���D� $	K�9�A,���������N�Ԛ���L��s��[���``�{�!�������\�M����풶�!Τ�L}����~��x+��jF��J#�����%�l�<z#o��d� *z���v������5*�5mչ�c.6�
ȅ�T� ;W�lpɜ�A�В¦0,7����V��������k<p��;%�����f�|W-U�h�-Q���e�FU��r�pC��)���WI���U6>߄H~�_#��	mTk�y�r��B^l��z�i���.�πU=�8���S�kq��kIn�JՒ�ɬ���sg�Ϭے�]�E3x�����,�U��?4�>D���,A孳W�|�f#cP �fM�.�����V���(b�]Ӓ./����ME/�V-��7���2fjP��2��KlZN��7�Ɏi9�8�yӮ�j��n�yHE�#Okr����p�X��z=�$VXV��"L�~�
�Qf��u��!�6�����dr�0�^]��.t������GŬ���, Ĩ��mCV�k�;�`.A?KF�.�*��~�'Pm2>eDJ�RA��V6c+̦���t�Wf�~)��ۮ$��f�ۥ�KȽ��b���Q���o���O9J5Ź��\}<N+�h=Ύ;���(W{�킕��#�;EA�1���hk�54TE|�ŴRԌ��*����!��	��� �S
�s"�y(����"D�V�#v���W�N��aΌ#&r��3��D_2t|���4�l���b��53L}��;��#Q �%��wO��O�����&�!D�1g��DT�2�B�E@ a��'<e8��~3���o�uL��d;�B��Ъ���F�cO����Z�)а?-�r�խ5:ǰ�澁�kR�4Qbw��9��!��Di�����gY�����������f�����Z��ux7�(R��}
l3_<������g;S�o�ue�N�8S�~��$pд�#��w�{�R�D�-6)(^mܺpaj�Im�a��fE|+�#�V�g�js����-@M�Pm	�x�ܥe�V�ej���0ϸxb�i�,Z7����y�.���|�,�wvB$CԸx������-�)�b��פ*)�~��T��g���T����&���ӗN�p�Va�0݋�j���g\��c�X��z�c5z��IH"N]�!��q�џWG%�{�)��ǿ~E;��{'hB�=�9�\�0�Hf����:'h���}�$�Z0��.���i8Q*�N�'��;���?z����nC���H�*(�� ��̌��}�ѯ0����)K�B"b��F�#D���ud�}�0ё]�+7�g(�:l�M-G���z�@�߇+9��b]v$3@�}%3�?¨�z]%k���c���W�Ƹ��	W��mQZ+)��2��_�ϙ%�����1�F���b�%#V:,�"��A�[b@���2d�U�2��ImÏ�	j#)��`:E����A}�Dy]��F����+��q9����U'�X� �5.� ��u��"����M�5a4jJ�G%8��6���H�h�Q��1���@_��(%��F��[#�Zؑӄu4V8�%u_��<�p~.ϛb�����P׷����РQ�n�U/�n�	��(|�����������$��y����6=���3�_A)��NH|���^�d����AV�� J��2��y���1OR]ξMuSU����1�Ǒ>��Qs�}r�q�Ƅ���:@K|��� .��E!����;kգil[�\��d�G�g���d�OM�.�ON4xܷ�}p�0��~\K}#`��-�;�\m�ƥ�����4ǃ�.9��h��@�qִy ��D��*<�H��`�3���4�3I��_k�R��`�h�4lP1����]�ԃ
�Ҧ	·j�c�~�o^��t� �h�SR�<�Y��X�/!����G����U��ld�:���������>�T���A��zu�r>�y��o�Q?��\_2��M�z~^� �p����̤L8%��1������n��	&�E��h�� ƹ<(���g�-��A����4�j�"c�����)��m��l�V�<�n%h|`�����,��HB`��QM�V����h;Z΍�A�7C� �T+X��n=���E�]���T��a��0&dQ"_2���T�Y2z�ضZ������d�Ә��^P��c���hf:�<����Sӎ�ވC ����,�V�	��|���d�a��Y br^�F��i����wpſ��x���R3]��:"1!������y�	JE��>�UB�!n�LxM�RTVi/Й�UV�$�[.լ���vT�@��N�m������dr*߇�	Y'���Y�9}��P�uM���ܰ�C��c�G���i�ai��Dj|����	���3�ݤ�S��P<s�����gf�`v�m����ϑx�������ٍ�5�� ���K�J�Jm��&i5׈E�Zsa�8��2ë�Η�#�����Qg9�>�(�m$��Y���#:���� �C"$+bȞ��
��iD2
��@o{̤f����/ ����Bf#�bM�` "��3�I8�%a�%�t&� ���g�ƯX��6�&O<�P�����!a�`�_����;�BHjs9Yo�u�)�{T���v٭P���g��t��㏳��b�T��⏨��w+�W\�3VB�38Ӳmx$���Z]{Z�PZ��P��.9Ln
�|En�7`9;�>��wנ�7�h��܍kN��(u����JfA����Ȟ���ӂw;9}�8oK�B�עor0"�O5ㄹ����tOW���Ǭ�J~/�)���:��'e��ׂd���L�Ӂ�6�K^�T�����.���:%���j}��h��jkAg"9�����Ϙ�g�gN�3)l��-�����~�aN��Ͻ�Cl�h��=cGa��h�s�!&bc�"Y�C	wRW5�7ɫ���d�;R`k^�>�bV�)G�� q��	�#
��u���R�L[�{���r�-V�91Os�'bhY1�Cz�-]����������*ʀ��_�T�{����+� �Ր++Gd�� =즡"��-�R3���t%���<���U��d��R���D��lMewe�U��t:$\%��O2�Yd��r!��u�^���H�jPus�����!�N���*�����]7�}K�����3�+��I��㮅��e�×*����
M�i5D�|��5;P��
5�P�R�elh�޽����0�C���?{��5_�¢m�ŎC�v��0!~-�6�3>:��r|��N��^�@���(�Jj�v�B�\���kB�����u���r%�+�#��7w*�-97���yل��6#T�c@iҞ�v5��є�!�Q��q2��p�b"@K�Z� :��V��T�gD��S�����mlW�3�M�vt���rʩ��t~�榘�4�B����7ƕ�Kr��"On�(̪�R��\�+��`ƛ&��2�[0�u�|�;����<n��I�v�q�Q��*#A��I�S�ڿ7�:��r #��U�aY�;;T@pط8��*ґ�e��*�R;���t�8�C`������� ��Z���Z�H)�@Q9ib����0���Ԯ&�Y�+�/�]u���S���H'"�SUc�^z /���s��̌ʁ9g!}F���q�z��<��b�EU�|cq���g#SƢ�I��%*Ⴞؼ��;����M>S����2��N?j`Ak��Ĵ�׆����2�uw��5F,q�R��bͱ��_�D�F@%��0�[P1�M����1{{P�Mg�!S�8�Ud�J��Stp�R��6�����m���m.����^#���1lXj>�I����I�"6��.�jE8�fo�.煎�<�:��[�$���Z��j95����V�H�#TfQ+��]b�(�E��x�F�)�w5	�u�u�8ұvpݴJ]V���1��9�k�Ut%�Ω��',������T9�E4���JVB���I`�;����΍±��a���\d�հ��pJ=�wU8��FJ��s��-_��oV����F=��7��s�sꮁB�U��t9�Ҭp!Ǽ(��
B1;~�c1"�1v�L��a �8��E�JME��q���?P�	�'�7�L��pͯ&��1���5�~�2v˅C��+� �`4�E�r�� �Z�ps����k�����=N\�ܹc#Uq#�ӗ��0��4�ncn)MH��t�~;,�[����3n��
�97�ia��5��*Vn@ {D�:�:�8u.�~9�2�mR�U�����+�a�Ŭ8-�
E^'ӝ]��()� �|��x瀺,�	�q���޴��ꓤ�lH<V��F�&���$��I"�qQ���R��FBØ�y�V�oO:6VŻ�[X�ꥦ;GH�������I� Ob�x�m�]�,e�@R6�ò�zM`L��^���@Um�.���_k�']I}���C�<6���R:���ùF
m�T!�o|F�)��U���g�Smu�S���Y����x��:� �j��TP2��5�܃i�
Ex�����7ڰ�֌͖3�6d���E�3�,N�q�o�I��77���c������6hzf�i��� 򍸯�GM#!y�S�/W0{�#OZt�S��u��Vp���s�DcIs�M4v�B;�h���B�f���w���@�_e���s�~�����np�P���J�LYkۿ}E�:S���O����MF�ynZz��+�}���L� d����^�<-'�L����cU�R����`��?�NW_��c��*�����?9�)H�1��	�S�]/��ckJt�I(b�L(Z(.�a1��eXZ��AR��Q�a߃��� �q��!+jm��w��Uv�A��vpE��Q= �GV����ξ6�%�6�D1���C&�AN����hÖ�iF�?6�q�B��=S�]X��?L�?�X��%��;���~,�׃��ۙ*���+1E��>�K��u`��i��2Z���	�:^��z�_�W5�m I��iZ��Ln&�N�/c���y� ��ƀ��WS�3��
&�f#�"�%�o3H:s9ѿ͢K`k�E�ny~�{#����7O�=��x&-����b~2s��4Sr��+BA�l1Sv�(���IW,��}!(i(S�ɬEeG/��B����Ұ���op�_�T՛�w��� ��}����ے��%�+8í��ֲY�]�=�����G�ݝ��fז*4TB�6��rM��*3h��n�4���']>�A��0�	�7
 =r�*l�����V�%KzD��[hp`�B*J��S���;`����6��Ӣ z��s*���I7�i|#9�I�6w����6�u���o��!�Jά7�6��m�sVA�y�S�"�ts��;v��7ǻC�嫍H���ێٛ�^~��F ��k����r����p�$N��}�KjUh�{~��8s�&�배��Z�i�:�)��ߡo����um�]�sQ��&$oSd7�PdR17�DF��_�p��cPCf��lĿ���h�{7�U���Ý�?���G�z��6�3O΅z���zX�1�w7��<��m�zz�@�.�[�"T��h.�G�f�)]�
�GA��N���Τ/���M��:IEm����6��[� p,�4������U:k�*M!��C��
�7vT�}��[��_�@ʚ�O���`r��(� ��5�^��睹��:����L��kx��l�i�8u7lؔ�,�� J�� l�j��k�����0f&�[6��0��|�}��2D#����H;It���b��lM����Ʊ��泴ޯ��1p�؄J�aL�]|S�3 uo�n�9m� O��Z�3��S~¬�L˔��S
!/R��!<F�k��e���$rS�M�z�.W�'�ـ�˞t�j^�v�yd��/��>y��/�38NS�	�����c��a@�0�r�]@ҩ4e5��O��_i�Hu��������,���k�^6Z���\[��P�Mz� �z�P��Y�Q���,�9�q�i[����̸���Ͽ�:��,�����+b�M�6�["�5�?��%��������Q�:4ͅ|��*�#[gn���#f�H$X��h��"��V8@z�Fm3@�m����-p|��J��;\8�b�ZA��~u��ˆ���������eo*�.�Y#J�B�an:���;��K�a,VBH��i���2#�Ĝ����� ��4��dQJk��%FJ���S�$*=��Ư�Gn[8�ǌfOj�.s?S4��ϕ�G�_��vY7_T�^lA�eYѨoDn�=�� �X��	Ti�{��z��0��Ee�J�e�=$ܣ���ݑ�$~΄�:����,ᐻGxk�쒼�͓ :!��r��<�~��CcV�6����)|���!��[����W�or6��2�=�;����agWJ��F�h[ӆ+���ɘ�=�<#ʐՁ�"�ޞqּ�hv�V����"+nV�)-�ƚǣ=�Q�����:y�?�l�:')����+�uOV�K��}��ٍG�k=r��mC�R"�+�\�lC�_��_�ν��������W�/c׌?�w,�]�:�/~6���n����7v�t-�H��.�-�"N�{O=�2�Bi��Fu��
M��٧LJ��S�d}��:��쀰�(�z�Ln�&���:��-��H���c'���'U�ycD�n{��,����Yj��¿�N�ʶ�U��	uɨ��6U�f��8X�r䱙X����0\��4�("���_��X*%����:�{p�>�Wb�V�88�����iP��.ɲW"��,ҋ5ȬJ9����p��óțV��"�m~�� �']_3���+�m:5��@���`p�whmל��P�ԳN94~��al0)��y�)#��TE.YP���z�%<���F-P@aI�W��ͨ9`��Щ��m}���^霡��&U���J�S�ERP��PԿk]���>����6�~�SVx{AyQ�ܿ|��~���i�G����l_������fz�\w0q�)��4��"��6�~>w}G��4x��'�?�nMY��頫W�}/��.�G�D�-|�����vt5RI�̰�.��U�#�9xz>�带5�u8�ԶS�H^���
��?>+zD�V��,���ݔ����ݳ3f�V�I+^`;v�q���Җ]i"_��PxZ�ǟ���<�?�2��#x�w��P�2Ii�p޷��B�2�jIp��Dj��?�;a���ˢ��V��.>1>���wD;�}�6j&F�-��"�4��_������鷥�����L8���C.#��SWC���+CyHs �2�/�z:���6�t|w[ �.�j姊^c��M��>����T��]4�La��!�q*��tbZ/I�_���ύ�>1`ȓE�3K�Z�5+��%���#�&���s{(��4�(�������'�To�����(��!g�ߘa�94��X/?v�8��9Y\#��A$�8�!��:���pc���y[���ᰥ.yG���l#�lt���V�ֳD������8qOސ[�ӱ)�!1���,��U���9_�u��4W�n��]����Q�t	gŀ�Ǵ$l���S�FL�*�	���%\���Z6엃C�:+v��!�4�#\FR�q@��ܠ��?8���9D���=2l�D���ޢ4 /�C0�t�a�_~'��:��W	�,+��������F�E��<	%��t��Gc����>X ���^�/��R�p�	�O+�}���rk��H	�`�0�U�
�M ���pOj���Y�g��4V�:[�0\AӡH���e��W���Zg4ݢ�?������窴(e��f��s��\�0 �1�_��J�H��/�(�jb��ݽe[r��|��ʔ{�ЀG	�\�p}=�6r�O�1֓2@㈄˓I�7=HR>1�1g[�NW/�)��G@��h��}�ōK�e*ڂ>��8I���,�
�FD^7�2_7I� ��>��J�/�#T����R���|��5�@��q�o�����|,z�%�ۛs>~>o;��+��07IV�\ (ܥ�L��<�^_�R��8��١)wqA��Z?L�1���)œ%J�2�2P�|'1B�?����p�o�L"��<~+R8pu� ����-���j�&`�f��`��>அ?N&�V�A��=��'E9�c��73wҽK�vb����dL��5퀠�f���͆��ҮKG9U8�O������;ee���bӅsY���s��_�OK<n�_�n���f�G����7��7��@�S�R�Ed3P(�7�"��K�S����
��|�v��eo?�H;@�F�.�q՜�c���Ѫ�v� ;{���Q ����Ʒe��ŧ�c]���OTh]�a�]�CAC���Gwb�$iY2Q"�{=��,O�5��skG�F�G1�B��
�t��9���|0�8��*ŉ�u��h�b^�.���G�}6¬���$�'��aZ|t;AMQak2����d�'ߐ��ڸ;uUT;��<����p�߽>����q�v�^���@RJb��W��T:�(�/�{�Li�[���a8��޼v͂k�[Ro6�v~؃ʎ��}�˖�����a�m�u�E9{F� ���M��\H��Э�~7K`}	�	U�;'YsoS���� b���E�@OZ�HB����3?���A��U�0�������Z��γ#���@���^�Y5�Z�ܴ%Y�)�F�����I�L�+�Fsզ��,��e>z�$�I�=�^R�)P�S��g&�"��kc��.�o�x�{bC��������s�Ӄ5\yZ�)�YQ7LY�Y��~M��:�]�l�1��U��T�! Q�S���.)��.�76�l�bs�G��"��)Z��)x�u���h������巘�J�gU��kd�r���`os�iX�0��4�o׿�*�ț\^>	���i-Dڌ< +IT%��^?1��q�5����0���/�g�_�X٪|�RG��n�}Z�"VN���n�N;�~P/�k.+;Vh=�k�"z�|��x�Fk�t����Í�h_�:l�e�t�X{���*�Y:�T2���\�9q����ܴWɼ��C�U[��I{3�KH�J,C��؜��*�G �P�&��j����1Z��/9 icw=�����9I���{Gy�+��u ����d�NgX!� ]�y�a7��@U����PR�>�dã��bl�\��_��
���{��0��n�b	��xv��� �����`���j} �u_lE{k�U	4��1���#��hԍN}�V��$�-�<�f�{4��p):���������.O��(�Yڒ�t:�G,CE,򫩠2�A���]��M��Rc.3V�pA���O��j�)�����O1���؊���/��hc-���sS�ƻφ>F�U�6�q��� X0ș��0��?�F�V@)����ި|�,�S��ȖI�S\^����h�wf0\qo-�P����8�^ xZX�,:4:!�Cw㷴 竎���2g_=s����,֠����pn�5�*���xQ�Q��D�)c���p���R_V�|�VZ�	�bugB��ݷxָh����Z~;w	\"�:Pz1q�7�?��m�?8��p�  t/�B����b*��tȔ�	�|���@�t�Q e�U�^I-۾�I���v��&b�f<~�55����9����?'�س�1�������}�||��E�)�(|A���ow@r�g�}�o��`I���4T?��u.ғ��Y��h�=���
Ρ�uM2l�iHxR���T(���B�Ƥ �ZX
��2�j����C^�@�$}��>�g���<ŕ��]~�`��݋��[	E��j�� z p]��������\���-M4�U�F"�?]3ʢ�%��z��7?^�=�d$�¢+Kfdu=�H�KZ����mJ�m����!��$li�r��O��U`�huBfd0b�p�6�G�eH�e��;H�E^�}� d�O��<�(V��K;��:�G)��*���Lp�2����C�#���oR4�ib�9׮�6��R�~�׻k�uqA���F�R�����^�4k�?C�sѥb&���{[�ׇ4}ϛ5���ĸ���r�������σ�u�c*�?��A���H憬@�/�U���#�}�1q�օJ������l�1�">��]c/_���zz���W
�(l+
L_)�=^	���S���@&;wV���-����=uX�m-n�)_i}Mi�?�Z���ε��W�"_�9Fy�;9�3��+�-�ȾkmQ�ˤS�;}�ыZ�����b�g�,:M��{ʤ�P���y�?e�lc�0i!5rE�����^����=��l�ސ/�ͺ���r���U�]8�!�
��B��H+�C��c��X	@�cK�P7v��|Go�m%f�L@���6�`73I�މ�\m���ul�P�-���>n�V��8���
�o[�u,o�ޯ�[|п��?@��ORvt������x���ZI*`k�:���II��Q����k��$��kZ�l4���:c���~�DN�8>�/nt���4!8S�~��+��}����T�2����&ߗ�5�o \,�0���H-A���yc�1]�5�c��޳
���̻�~L:�r:b�7�+ڀ�N���d�:>���[��1F#�!f*`˞0�$^���}D�� ���+���CC�̴�� %��yWWz(�y��WQy^�(m:�e�9e_�z��L{3� �y�x	�Lx0"`���BG��=o�'�q`[I��D5ip��N5xO�j�Nޔ;���zX���IO5ɲ\�l��U{�������-�W��kH�Iv�;�	r�TU�%�	�ִ��J������9�ʸ�M�,�ֻ!fWѐLc��ܮiꜣ��r�x� ē^|��g<Ķ� LN�gR��ʫ%Eѫ$žtl�Vܭ��+��<��۔�Id梗3��`�ͳ�Ã\?��!��p��|
'�?ю_h�
@�d����a�EȆ{�r|�pOA�&��"�y�����TR����;�ˬ]%���� C�`��#ѳP櫲�Z��Y�M^�Iߝ��a��$*�C23A���H}J{�9 ��ћ&eA�3S�v�E7{,�
�B�$z�I$}���D�`2��+�M�ed�@r쉢+��<D8H]r��ف�pw�=�-�Z������f�+d�����}�	�Eƥ�cK��q]�������w�^؀�Mx��0��v7��C֌vG~벪���Ҵ�2��^\sO����1\w+����L�d��`�P����;��	����"�^0���A&_;R���6ʯI�[=b���'Il�,K�҆?�!*ԩ�矤���%x�O�遼4�,7�7�;���ީ�ϟ��G�hP�5�3A����Dy����ű��Vt����n���61:�ҟ�R�� ���F��1Raq0�ۅ����πc��n��z&����؏_͘�ζZwdl���@�$Ӊ�]gl��"����"Ke�o����4��Xa�JŦ��ҫ0�?J�⡻_4�l}S��u�
l�ov��VDʌqBЊ;t`@����Z9�L��a�fA��}LZj5����XR3'�g�z���-@�߽���p�қb���������8�fgm�яi�c�|��!��v��^=�b��VvtzM����`C(mCV��dxb���P
�@�h�șW-�j1y ���X���&����Z����3�/T�͌�0��y5U4U��d���fA��E�`C����ŵO��HY��iB�4�È����j�j[T:<����.�[��џ�M��=��h%�x%���~ �!�
�܈����%g�����l����c�k*ibGQ��dT���;sh+q�d@yTa=����0��s}�~vի@M�� d^�ٕġ+��{N0���SއI��2|�D4aR�;�)��<�̏4J.��DV��U�VM˯�M�XHV_ƚ#G~�XO��]�FU�A�4�m"���P	ZҌq�1fj,RMk=��I�@���a��`��Ȋ�	�� l)�C����
��O��	e�R�?��
��g��1�3+�`J��D�ؼ�� )��%5��P
�ȄV�%��yJ:�<ޞ>���*э�]@����&����J]�|\�b�x���C��|S䁎��i@�������"7F���6z�vM�7�=��Q��K����c�C�p�_Ǒ�Ŭ� ��p�������5VM�BV�!@S��_��qTu�Z� o_���{��pA�8��步��&��[��{o��G���5ɣ��a)�!�^���сĎ���x����Ͱ3�P���|/������,��Vp���B�F�^�Rޜ��0�ʚ��'=�P�t��m����T���v��1*�����b�*���i�����1G��Ӧ_Tm�z�/6�oG�+�z~D�����ye`��	l�S�v��ɋ���Pv�jUأ�ٹ��ҧ����P-��t�xߤw��>�]����L�xrA�vv��W.�jy_���O��A���-A�5�E)����I��0	+�|�1��v�$]�m.��@�,릉#Rt�H"Z4�!���k,���X��ٯl嗓Zz�⥗��I�k.�4����Gl0r���)t��~7c����]�%v��A��юKJXo����1@g(�[��v����qй���g0�V�����/���|�*R��qT�H�|�����ӊ��-�s��uɥ�s"�$�pg�ƫ��y�ND� �Kܩ2����<�uX�޺^Z�!��f+H.&��ئcq�
��ܼ�X݄���&"�p�4�����O�8E~�����>k�2��(h5"�׿�xu�8@ �k"����*jtu�����$���}у}J����W>�ڹ|<8 �h�83�j��$�@Į!U����-�>V�L�)�����{�+T��A7���o4������ ��F@m�
��[�V��+����]�7g(�Ψ��;"�>"AоP�ꝶ
?X�W�F��|�>��D���ʺ�&I)\4��q�N�TҚ�r[(�����ԇ:�S
Ex���	N˔t��	�Β�f�{��c�" �D�ܑ�}7Qa�B�qkeD���܅�B���h�E�L��6��BxƷ�۠��9��l���������$�Ƴë���A��&�y���0#�v*�cfT}��҄��I5�炱f�4��oz�\/qnٸa��l5�gg�!J���iA���@��6�7���"�؀��sf(��n���^d���]��	����Y#�e��ij�|p�Ņ�����7�'��a�mI���G��@��̢?�x��r6�/(�e��of
���*�~{.ey("�@T�#�>������@�v:�lKV�Q�9�&�_���H��s�-���: �H����H736Zvf#{�P�6U�K���T�PG���hb�u�wģ@�`�]����p~��iC�-(?��.���o���,/E��<z#�[��Q:�B�cp�t�N�	���PB=���rl�'���������>��yY	!6�<��^��i�|��8���ْ�҂�J>��E_�}�0�0�~\H����E�h&��T���I��Ѣ;���}�>9k	�O:ѵ�/q�u9_ʮ�6���|p�
��1�Y��p��/�9��3�=`���͗b� �x�L,D����ی�~{&�!��GF��2y�5fV�N��zT���
)͆�Ʃ���6�X<�L�HJ��V�{ioe1A�\N;��1��w��X)Y�d<D[J�������jDK c��6��nq�������Űh}����Yg�*,�B�(p��Nwus�[cǞTX�:���h$��O�pkFy�a*R�`���R��n�	��Qw�~�̈́
W 
�|�d�/�XG�~i��Q^���^�?H]��Y�KX�'�?�$�ga~'�n1�Mo�2������DPw6�ee�4�G2�
���{�+���W��\1	,�_��S�I�:�Jm~f��'xM�(
�aV���Z�g@��A��|�q�(V���7�0�p(�hc��WR��>!i�1T�#�5��@�K��g6���A�����|�3��S'jd`�����<3��d;#U6��(b:���8'��Cf���&C
~i�j��H$�
�JvO=W���l
naI����޻�PK��T�����^qI�KS��'+��Z��%?��*׾�y_�x1hspT�=Zח��u3C���=6/�}���W��:}*,��Κ1=%~��=�+�=�o������LL���Q{��d9�b�$�U��C�����.ꟊ�zƱ�.��hg{��k�oʦ[C�$�%��Bu%�!n�f����6�o<���b�?�R����lN�5c�*�>z�<�`"j���%�c�0��`�iS���x$Jt������e�SD)�����]��Re�A,@}2w� �����
��91�DVHi��h~n�CSė���Ft��c�����D����ǚ��,o�h:��$j��阡7�H��y��z��7�i�X��W���Bt��Z������ 	�5K�=������ 6f�e���l���nS����+�I8�#�8���Yf��W�i *^b��2�r�;G+J�`����7���geej��D͗��� y�
т��y6w6��p����B�
m�ILt���y��b�V��jUL��Ϙ�;ԃ~�>�Xc�B����Ҭ/�tw.O�]�ƛ������j�kG%�������Ј"�Z�i��r�B����%�w_����Ze&p~�����L���Hb���Q�a���%�J��Ʈ���X8��aS�?>�np���]���?��Ll���h��`������X9V�h��}���F��]�#�mI��ݥFWJX3�xB�&��C���!c�w�ţ߰���Y�)H@9ՠ6�$FK2v��V��ۧ��i���U�WV��X��Ծj���p���k�%�I,��hQ���X�ً,���~�Sy��G���\��Nm�{e�ʵ��W4WJZ՛�CS$Z����KD�#?)'���~Ǌ�wݐ���ջd�3��M�V��Ư�I�����l��'X���& 9R$�"1�%��_��Hk���" ��懒�)^��^6\�e�+�1��CV��³�ⶖ�= �m�$�D0�U����$�㹺:�\�i(Z�������U<S�������jh&���[C�D�VL��R��YO3	�r=��#���ie�����̊7 �l��	��8�m�����d��2kْP���[���%�,L��
t�)"�0����h/�t�O*w�n�"twl?i�_�(*�o��1sF���_aV��0�ѱ���]'~�nF�$@�����=�8F��m��&�͝'_:7��D`Ҝߍ۟_<ڑne JY�"��~`pu5Z�-���g��R�4a�ּ�f���hE�����o�~m�z9�xR6,��ʗ<���H�[ms�v��8jzF�R��:Z�#�z�߼x��8�ORV��N�/�S5N�܊�9F��������v|~�1�����%|��Q�J�PMmxm{�5�0n
���Q�\�+a��8�u�#�����]�N�nȪ����ߛ��@)�)}���I��%y���.�����z��+A��;�������LO�� ��M��S��Ѐ��Ȕ�A%�&��Ein���+ ����\H�r�>�������׃%_�Q<�~�.�A�SN$��O��o��'C�|=nf���!`](�W���Is	ap�9-4����"+��KPY}Ĳ@sB���w��JL�q����5�_�����t�=��� Y} gp�v}9'MZ��Bd��-89Q((=T��1��X�PzK$f%��1�^Eu��F{����	��M����goLoS����+f�I���µ��$�=���r�"��X}�#��2�F�4����L�~�	�cKrW@�!����k:/��J�[.1�l�cA���w����<�}3�{��v��4Y1���1FX�����n.�8 +DC&K2L�>��YBR�7*;nG �%���7�W�\��ܮ �aP4Rs�@�<��R�<2*�%Y�pi>)�,Bl��w'��ppFY6�b��H� �f@��y�y��X�L'�����a�_S��R��ƃv�T%Dw[��.�e�i�T��|����}K�~�ۗ$�4���:�����Jr��3��01���������l��y&�%8�݀�\+��}�T#�&�̰���Xt������W�˅��3�-%J�~]���R���0�Z~�>=70H��R�x-R�9t}
wQ}�*}*!��Z((��T�R)��DH�h�'0]�]����	��?~���`��"zR���[�����	Ͽ/� g-	���9�;P��c�]|�N���}�1��w4��6�d��
-'qTTm䥦Zdk2�����

�,���0r>���:�����Ϸ+�Pu��GǢ�0�?`=��	0 `FV��Ӂ��!]f�B��9�ԟ�DSDFq3�4{W�/Z�_�a��tfr"��� a`�{�}�ȝ��<��F�4-�6��R���C�h��7\��[s�>Q��_�6�iaUes����"$�U��awڍ�ؓv�b�U^S	��[����W@1k��JmfV'�,�1+�	�Fm�ӍN�ڦ��!J��0G-s;��K�2�?���U��%�o#�jJ�V潠65[�l8U�,$?h�O�Gk��b-ҷ�����Hl����N \��������@6�A�8 e_+�J|���:�4V��=��3�av0�ϟ����5���W�.�,j^mM�[(�Y��?����4 �d_�z��7�7��Yh�e��:�*�)I�Z������RG��#��ʒ��[��L���n*D�iWŒ�����L�|4�����e����el�`���(�	�L�OM&a����bn>=dy�'��J��Wd�d����@q������t��s,�[�Ք�͵�W.}>j�n�����xs ��������(�buwv�ޞ�e�z���9�oڳ���+,�pz�zs,��8����@��ʩ�ҧ�9�Z��	_�!�c�<��ͫq��eJT���Y����� ����kq�ܬ�OI`'MF�p���1�Ϭܫg��u(og��B�uX�7�6�ڕ�f#��W��D���������§�컾�ͦuyu2���%��x�*�BI��b4�6L�!73���{I�w{�R�xPK"�/�#S�oQY��ÖTf�� ��=���-)s	Gpm�-�^vg���F��%uB��E�;R�R��`����h�sfz�D�\<���`���/�[7h�y�|.U/��M'�ɒ>�f�,(�г̡�F뤶�#��]�I�7*�d�=�of�������ouuq�T7�����L�3�ZTv��j.=�ʵE��h�@�4�r�|��d�$QfF�Ʌ�읝 lF�M70�L�w*�B/&Y�y��Q���G�L�߮�L+)��^��gj�f���$_˭��y�}���*��1u��E��>Q/�Ee��r�1��e's��m�m[�1`��J�c4a�X��ަ������)�]�ל���Z)��55���� �f��(����aZ�X�qnS�X]����<|�k0�⓽m�E'�Ẁ�Z�����up��:�U�d��feW`	���K��7x�v;@�!y���:�y�s_.gZs�^�I~�t�g/�s�j������e�wlM�oC��n ^���wuY�������غ��+�%/Iӄ�}~���8���5V�;}i���HW�>Myez����A����V�(�2�2(��.Q�1�ʚY�whd��K!>�I�*4@��1�R77%��œ�T�y�3�Ө���h��؈��D��'(��k�-�.�{$  ��mt=�4B{(�$�I�9�A�[�e�����Y���J��np����e�`�l�ц]�f��ζ6���ZF��Qv�u�X�zz�^��|Ō�Y��'�U���������<zƄF��̆x����ZBQ�˄�ȘP2�Mm���o���*���{� 1s�GY�� /,��te�V����̜�ѹ-'Q��>!��~�.Da��J@�Z�1�5�M*���/UC������VQ�����>�o%'��3���s[�7P����<X�Hr����U\��A.����h؝ǭv��d}k�) ���9�I$���X�B��-����&G'�9���*F���o.D3�qd�7�X������f/N�C=�A�y����ę
�<rX����Q7�eS$����[����Ϙڒ��|́6����3�N-zr�KDj=*�����m����41�E���
�o��7�*}ǲO`�������Ӛ[�kv%�0�1ʸm�<��r��×��@!g�F��(_F~���Ǎe�v�6�	U�Se��ʭ'��>�:��ue�.��ZɅ�T�\�]4�$��U�G�`������a��dj���o���Db$ã���R���1��4���4?)��IFwp���%\	�Lj12��o(e�)'f�#�V����E3�7��[�j�Z]oOC�9(��#�7hx@����ewF�-�}��X��սV_�-#�R�wrӥ�e]���6i�Z�Nx�i��5��^%��t�f	m�n�fҴT�U2LO�t@�����n$������} ̣�Zϣ��U���s�K�@	"��=9�᤾`���;8�G�Zp�y��_WaƆ�.�-��\W��M�L�<�G�[UM�un�2��W9]bdAW��vT�@c��ʉ���߱b������T?5'di�I���%��ɩ� �R|�J�W�HA�[�;a/e��A[ݲ�_���2��@+(|�E5R�k����LcO�6�f��ϚKJy�Vs�ӗJ�r�	ͯS]��$կ-��O��Ƃ$�ʺȶ	�y8����GDy�>_��T�A-C����Ȕt4����	�9z���'�z�r�fVX�
�׮�;�K�P6�²dP}!�p�7��������:@ ��}��������&s ����=�fS\MA����x�~��J�����y@�~�������Q��!�`���[�>>�S�
 ��G[�̦"|<��XJd������#$��D���G�	�4�TgC��x�7�STI���R�	6�r���ڎ�Nr��
N��v����-5�Q�RZ>��t�����(g�j|~W�h�D�\�1 3�r�^���� yͬ��d �h�^ZpH�*�#�-���)3���.Tc�zÔ5�7��cu!�8=��i�,�`f?��L��q����6��2��J���3��0@Ne��D5owvD
�F��%�F�:��2��ШTA�����c�#mq��m�MU���!�#hY1��Ի*�:�9�u�и�ϱ4L��JY��Q�̍��:yP96�^���Cjk��� ��ѯo��᭑��)����W�ъ�|�yH@Xx����Ș��;����qs�V����]�tLS*:@5�i0�ZKg� ����2�Cw铐�~���@�)���� '�#��I�gK!���9	�p15�ŤO��	8��F	��?��N�q��;��@ەl��G�P�o���Ҹ���Xg�C���ZK���"���x�Q�m�;��j-�1���G��?������'ld�28���Z[��P��8-�l�K��MI��JGQ����O�9ف���*qU���󤎄/o;6���>կ�v��S+��`iT� �n�y²�j��bl ��+A ����{fjk��{QJ`2	�˭0�!$q�V���P@����}!$C�&�\#1P@���#�M���8�ߤod���������ȵ�$�&O=?~�~W ���eM�xH�yc��T\�G9������A-��Ӹ��|��idO� ����8�X�@i*��.	�%�D��(q�|P@5&�	B`�d������(������[�YK׈����e�s{�u4��%����ߨS��ǍZ�a�����>�Ҙ<l�x�t�t�N��:�|4#�/,e�����\9H �]MƐ:=�|�}6>�Tk�\X9$\" �w������t�$c�	J#7���며ֱx��C�ƔE�u��	T/���e�#���rt>6>#���O�iP[0c_N}�r<+��aF���G$��Љ����zHV����	��^wD���"�Ư (��W���z��aZ��l�����A�x���J�C�=)��^ιX�/�n�0�����о���Ix�΁o�&�ɱ�3�$�H�αZ�A�2P-�s@J���	���(
�n�ng7��6o���%H��9(�Ü?�j��6��f�)�]�v�l���×Q8���j�Q|�4����>����5�L�g��uț�Hx* �'�j2l��#�1X���|�;��s.jAJ��ZEq@o���_I�����&r�y#�(q:t�=��h�:�9J���+Mέ`��N��������8�Rk���LEv4|�)���>�p�-(xAK�5۩ ͮ�?�&�o����"	v�?+������*���3Q�c�DQV�a=fh��jEe�s���n&o
��7�M����7Y �ʹ��{R.���)��<p�/|���t������7\�,����;Y/|���Sd�Q�x]���(�_*��.�BB����P^��+WM����c�Y�!�������6�@���������5Ljcٔ�x)�����L9�+	f|�߼A���k��/����r����r�]&����%�g�&me_R�/�b9I�P^�*�n�q_Ў"|����壼�����=;��H�$8��g��Q�b�]5방�7�e�P帆�R��S~����C�H��)z��4O߃D�b�?!X��F�B.T/�X��&��{v�:V�>&�?�&�ݖ���,�4xJ`Ԭj�;� �b����.ڃ��A�%'���Kr:���تS�2bG�e>'d���˫p��g흠}Ƙ]F��͒pZ��m<��ڎ�_��SB�"���kO���!���2Ӑ�q��9�h�/�����#]�+� 8�U\fr��⍲�|-���R`}֮��D�UG�2�z-<ZS��/X�m�6|�l�ԎPe�G��Y�cjfɬ��7��f^��\�/Q�cՄ�z�%�'(�|�'h[� 9�h�۲��}�|ѩzj�`��T��~��&���\��}/! 5ղ�0Z����E�)#�;&
�Z6�N�b{�-겟vn�n�e����͖��Sc5��ߣ�P�}�O+݄JW���P� ��y3T�u��8�[��:_��>�7�fXL]e,x���.~p���c㒅���� �
��