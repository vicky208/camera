��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:���[�S��Ɖ8��1�W��f� ��OYli5p�"m����B�t�PlA��Аӽq9X��j`C\�m�(��]e*2�k�bǭ
���:�ިRB�Zy�no	K�Oݝ!w%0� �}>�t�U$���D4[GƆ���<���Q}�Vn�~�|��W���d�����X���f��rl8���M���iw��i�
鍭��r��632�uqB_>����lOq���/�@!�$����A�r����z�1	�##^z��F��ڋV׵�>�8v��QMQ�%G1���x��,ޭ���FY	d�|`��;KI��KcW���qb��n|��g��hF�Lq�����VL0I�_��-ݎ_���U�2�˗}�ŷ�~b�r�Ì�Ԡ�l�߿�2s} a�T������)�*L� �,���SFߴ���@b&��J��-�?�8��>Y��~>�x� ����j��>L�P�m�*L���emxfq�1p��������j\�X���Y57{J��v��G���E� 0\�� YY�k�>��hy�������r�^PWLDC��O|y�PӁٳx2E��!��Tq�ˍ���8��	�v;�%}�zS7��F�f��ݼ򇞷��g_��i��}}�����P���4�YipH-���Mg�]!��_H�M |�jU��wG�1s���I�0�n켥(�b*�^�Ŷy���'��}�m�q,��X��q�m(�o����ß12�T�i٢���4��~����(�s ������J�،B���o�s�r{�A��x#��'�9�(qA��?�+GD�2��^���ː��X�D~V;����j����%�m���ȴF;.���ψߦ"-%�f�2�Ҟ�&"��Sb�8�r��6�+�z�EL�ҿ�骥�4�0z&s��$��Sh�~1��f�>ݭqz����:*m��TO��ﯟTZ�Sg�hJ�X�1λAKy_���V��	�6R_)2�����:�D��`�e����J�Ξ��=C��G�d/�Y7r]q3~�C�E5���#�B�A�2�*�Y�EVD)Q�Q��ذ��z�"�=;���-��?�p����s\�)4�"
�u�Rl��������i5T��d��{+���:f:yIHdF���y�I��d@�c��	S�ս���"1�PS��	��F���ؓM̟Q��r�
 �L]���<��Mo�V�T0i�������w�6��S�M2/Ȱ?�U}+'dS�ų!Ƿ�����-D�@�TQ����-�fllYG���n���)�{��kþ)N J-�J��u��1���Ux����Gl�R�r�kQ�)mG$��C�x9�"����k>ޯF�U�܋��R��|�'��0�8�hri�ʔX�KUg|�HHn�絛���5*r[�ư��qNf���&̩�)��_�w�Ѥ��q�	��o:�>�'�/�����Y�lH�b������g"l[]�׎��ܜ��.�1��0F6���؟[�us:���ܢ�v�W�gS�I�����_���E�`J'�8�|#��=q�[��j,�!껡��3��N�G.<��Lm�����<����m��LWt�eӄ��� ̰�b��!EXm�\���y2o� >�9j\? ��c�G�@#�7=���J�IG��'��q_3���^_]>[,Q��o�Y�G��?~a��]��8����j���Z����n�p<�ڃR��I�=zٵRx�k�c�&�$��z��Ze�XE2C%�4�Ξ�����Wˑj-�w��^�zJ�(��]Y߯��9�;�`�Մ�F5afe\��x�|+O��G1��?�v��(��*�h�.�6�v�w���O�ϲ�e��PV�zu �=����LQo����b���s*ڃ�P�X�l�OMj.e�L���S{�4?��AF%Q��o�h�M,)s�'�_ ���+U�7~0t=`���v� �؃�W�<޴Ȳ��ƫ
U6�l�r��d��ڐz�c�I��&�s0�3i@-#��M)'�H��*����&�����A��d��=F����M%��
K,cU��nY�S��4I��vKV������t��$��z��d�6U>�S'E��)��
�-d޼�|ZO�g��:��w2k�O���50QO8 <>�-sG\���wׯLl����͒�[<)l�1�E��_+���Ë ,u> �|%f%J��ۨ8p��D�Z������Zb��9�	�p�>[���8@�/�a����Af�=�
n����7o����6� V�N�)�ڞ�%'@�Y-v)��kJ!����2�P�?{[$�_�7a	m�Z?������j!PW`���2��0�I�Ҧ�	��oݶY�����
B�����M/�Oa.�U�-R�I��'X\	 f�F�At��f,�*�'���d�߭�"���	巩�;��de3�������'���?lˀ{^����譾�Kh�B�fE�ߗ�DIj�M��~�(h�e�P�L%��(_�<oQ�Z�����=��/uQ�V]��a#�e��:�5�!*��Y���
y����%�H~���)����`�� t�Ş��Z%e���yx؀`F ~P6W��;!�A�VԊ�9S+`<�~�*`����xעV�5����\��2�Ǟ���5�f���M�e�('G��	�6��p�-/�ID�>Z�}�9��S���A�^G��Vh\\����Xd�4F9?�vSD3��
X���5�;6,#�ZKO��\o�	݁��xY��xv�����0�H��v���������V�o^:]z$���L\/�Z~����� �q֓��V���`s���5��H��ۄ����ovr��PF!ּ;�c����T�J&�ٓ�����&�Eހ�[�:�?��t�Iw7�#c�Rt���d�<dI]}��Uϡ�O�����D1XҏY���*f���X�u�7Fط'���.��A�R�)s�kO���+�<�P�� cw)�,�V��;KpSk�M��՜����Һ�{Ο�5�YB���w���,���թlʈ���H�+a}8�::r�>Y��+z˨�,B�����4�.�f�Gb`����IU�I[�X'��'mn�9�!oPd)����2�b	.���à�@�0��uk�/W�Y�/wd1�+e������*�c�2Sw|?�,`|4�b�/g�2U�c�� 2�K��d�0fG%�@��z����,#���')P���������H��
�W��gD�m�+Pp)�J���+#�iyw1馫�3��/ٳ3Z�m�����+��t܁��^��4��~)���.ևr��u��C�0���ML�k���:n���	�VP*DH7OCw<��	%��NO�s������F�������0{HE����������G}9o��������,QԊ�r6>�Z�"A�U"Gę��#gϥ��wr*���G��\.׽�|c�v���悟�!h�X�4$�N�:�m������./zA>�ܫ�q3z���z2����k��R�Q�p=�}?>�}�KS������5����1�}����G�_߰I�_� OYGWgs7��i!�W�sB	[�I�-�c ��NfDQ]�S��w����=~�����oמ'�O,�ه �7M?�`���1��gˊ��M����ЇN�KV��թ�e�����gU�7�O@���Z ��T��Wr,��QԔAI9��pk��\��G�<^�M�W��B�}�N�z渀s��߮hh�k�(M~!N-:z�����L�
�*"�#׿-�A�S��K�Z�RBR���
���M�.��-Z�����j���`�3�Z��X��L�L�S3X�F�6t���@�\D�2�}��&�c���$�Q��ש�m�n�O+�B�_����!�w|��!���Zp+DwC�oR�������x��6�y�x�� ���n�q�kF��&e��m�T��1µa:���Χ�겒��tm��7��-Y�H�.$
��o_�^�J��=Y��~j?#�E�?p��cqk���͢r�k� �CGC
B����wCOP����%��$`h+��$KdJ�p�9` ,�]�X�r$�b�c�x�ﺁ��ꓗ�x�m���Ǡ���4}X���y�T�I�j<Գc��`T���B�ȣ6B�ND�G����3���ލ�^����b@�]��W�|y� ��ˍn3]���^�p���=�u	{��' �7w�c��KY�� B�6yRi���M�A���ȯ^Y_ޠ�e��!�U�8�;N0t36�!H����K������MfJ��6��'��Ȁ�r*��������dM���Aޞ�����R��Zl�Y��5f�e-5P�v���6{㕗�(PepEy�~��bą߄�1^�JkD������`6�k���Vh�J쵒Ty��9����� c��W�s U�G���\���<"O���+�2m�B@C��s�>��z��+OƳ�0%)$�B�A�#�-�ֺޥ��kYww��c�P�~@���A��k�Ӈ��ښQ�����M
�qd���,�U�OX	�Z���2�A#
��^����1��o��P@_���|?����O���N��uĂ����[+).�鵭�`>��NED�����*��Zq�y�5�R���=7����&+~\�Wȕ��CU,-��F���̛I^=v��R�����tB��6W��|h��o`t�%�'R$o���T ���$�P�Ơz�����i(|&�K���<� �.9���K���Ci'&L�I�r-�0r9u�8�ƪr"|C�V5� L�b0�!&��k�?��,2��Ȇ[�s��#l-I�r"�\5<h���G(r��gfR�9t@=�(J��46��(��k^4�$��mt�Υ����w�c�#��+mѣ��`�z��M* W����`VeF�X`<��݈x��E��)��8��.�cFN
��[�:M�(0j���:���HN19�����Ԅ�-���h=�#@��{4Z��P��𖤷.��?�J�nF"]�6�&8?k��|�ɰ�I( ���o�$w�wtR�شH���������".�8�j"v͋T��M4!2˸16 x?�N�����Rʟ��5�P�J08٤�>3%����N�c9�~�j)�@��Є��z���}�`��4F��������Ɛ���s�@U�)�+�T|��t|eN]ye�H�EM�����⍱ܶ�)�|
�D���$�P��6���j��x[ٹvW�x���y��g�f�Iv�����w�K�p�������^|���WWptf����Y�?���1
#�c��mc���
_�,�Wj�Ә�P��^3�B�K��gY�w ����:��X�YC4E��/.v�ݵ�1�-'�����T+�_��r���0{��#�u4R�W�q��"���'�q�c����(r<M�H���b� �K��H�M�.�@�{��ʳ]�؄}r2�CS�*K_�eb��7��Ĳ�c�ʐ3�u���)�<��CKܭM�M�x����ݥ���ވ����ܿԘ]��"*Z�q7�i�[���yĂT^r�:K60I5H�W�f���vy|���"T����u�~��(�D���7}�Z���%�Ҹ�R\N�?$���'��'+�A�cQu]R�d����nfw��0č�\)��$�.>~�FjiK��uQ52�9������BN�5yq�����y�`����9œ����Z�%�����9堊�/tkX��5s��%��%T��^�G��Omx*^���_���w|�V9Cv����}����!z�!�K:3=HxjZ���o ��/ڥ2j�wʣ��9M�$T�c�K�Q�����hx�	���g�!*�H(M�0�s"�/��!ɜ�{0�"���ڀ��vR� &� v֑��3��hvB��ڻ�#4� �Cr���M6,�yޟ����4t�6��Q�g�X~Z�����T�T�Ä�J1�Xø`U��Wψ�l��`��{�F��/��_����qzb�@��4��bg�kg1��=��Ԙ��;5z��؛L]�u3P�X�i�_q���2&��x����8g�}B���OdXӥo4�zǃ�)b��EB�o!�:h�@/{��Ȳ���1�ICW���LXX$�L�� �6��i�l~�`^�)U���W����E��H��#��X���o��ߛ�0�g�-�wC�>�0�
 =�g��&@Ea��Qv�U?nUa�����m��~m�UW����=���~Z3Ȣ�a��Y���Z#�P��>#�.��:�0���+�Pe��bV/����L�nhS�Kd3Q��_`d��f�T>A �&O(��/΅R\-\d���O�;���͟�D���S�֔C$�(=ո��S@~%t_F�І.�4�{�E��U���6�����ƹQ������%Wr	ST�F����&k��r0��v6���`�qʷ��&��������5ģ�Ɵ����m�h=B�뤃�K��s%��{|۰8�N`�j�2|�����XC��;�*�? ����i�F�Ɯ%g�F�u�D[+C���E��5^S,�y� ��aZSJs#Q�4Ea[�!�]&�CSbu�4Aϧ"dT��9�4�8:����[ ��NL3�į�]GT[��F&�;v����i_೨Wsdn��� Po�mS� ������L��V�����*�w۾*=���B�R$gZ�,wS#��H�[�hW���C1\l�����3W�x��Ro��9l�.S`>��d�;�W�L��/g ��>�@s� ���4���W~���K��u;�K���@���l�M�)�ُ昛����*�����i��eK��8�-X�Z���M�-������p#�`�W�za�*�":�!s#\�����6��L��q-����|�>~�~V	����P�M��l�#�'���Dφ.�q?h�Nr<����M���\n�RK�G���x,��/�Z[��)���!
,��^`��#���f�&~���O�79����`�S�ڋ�ɤ/=���Q��o�{����G�:Q��S��� �=�G_Ǥ�P0 �;����E�,H�+�:��,ͅ���2U��G"��L�"[�7���X�?�|Y�t^���j�6��w�~��j՘߲y%�J�J��H�J��Y΄����.zQh��o��X����2���[(�"�ĺ]$E�e�나��/�ӎ��*�W$�x��w�P#��6���찿Z�+)����]���T MF���`�.r�y[���^�6`R���J�;�'v����D��
.�j�2P/��	:[x��2��VpH����P<Z}�u�Ol°
���(�2ߤӜ��]�Z҃���~Yӌmy��؜Bc�݀.�
�S�Zd�ף�2��>�_���9u9U�\e��&Ôi�,)���<�s�V�s���B���Z3�����N�����vk�3�c��U�}DX��R�]n��*������T�˷}��[��ݜ;DH�v�4�:�}�u�6��p[�טu���6���u~�!�܏Jt��4�e����5�F�*.��3�5L5Or$_P�����[��#4����o`X���0�A�:�~!$� �﷡���.�����EŔn��]��8�����h��\J=1+��O���R��T��=���fJ2���汫A��fC0����2v�U����cw�l�S�ϵ��%X���1iM�u��>M�$V�_�������i��א�uZ�2���B�2m�^��W���(�����Euk�	��=�>�kD{g�7�L����� �����&�tt���Y<�w�nZ�y0'Xդ��3�7��,Y�A:z��(�T�0�J�,�k��/Ҋ�����T����۔�"q����҃T��l"���̉���q��[QT�|�Ԣ�P*��� r���cƩ��X�]5�麀���>st���H�EͶ �Y�ݲ�Ng"�t�Y��>� �ޝ�0���ᇍ�:�wDY��%�8+�wy�b~c6��u�[瓚[zH�&�t���
�����Ē�m�(�/��Z8�A���?Hc�6�u�~
�C�S�&T9:�s{;z��.�ĺ�~��Eڕ,G7�VKo,"[Zn{��gV0��v�|��-�KÖ���A�����k����_������O�#r,]�
�"��b�'���9�`5�N܋;�^EAiz��O�MI�on�����EX��k�yKl	-[����.-�N��a����'��u�Q{��5ꆄ�+t@�B���8f_�v�3�Y"Ώ@��� ��&Va��mPCq���>1����,�Uf���N��e5��ڢwv��.�Xv�_�-�J%�b�V,�h�s9��𠽒��;.L3>��-%h���K�R�k�m�a�|��ד�{O	tO�S��s�Ir�G8"^�/�P5�j�,�.x.k�Fp��17�����2gQ����A��[Q:{���kmA��:��߂��w0ILggd�����i���m�M����4_\̑v��Z��Z��m�u<�q��w� ��i��a�C�#�'�#Xl= *�%���t�e^�#)19�0� ��&���pc��}؂6/�f��N��9���h��A*t9Y5ѳ�T�T� e|�� �~��ê
��p��-y
�AxX��/�i��>�2Gy����fx�-�e���c��	��D6{�t�2����/�����<�n#��!+a�����<y��뫬�hɖ��q����pi��o�����дae�v��ָ�|0�"��脾]'O0]��Olq�����m`*�G���f�&���ՊQ�o|*:��_&買����+�Ѱ�!8��|[�Ch�$��K��4�dy�s@�62?ߞ�6�!�A�}yGec):һ���A� ��J%��J�U�w�K��vj����3�>EZL�HX�x�I��vH�N�6�����U�2_�~Rf1��b_R���4���5L<�"��TA��"����r���w��Io�Gq4��;��&�*�{D�y�Ço��l T�I1�aiw��B|-5K�y^,P1VKO
�9~�m�2Hl��@�a��I���U8Jeąh�6���I���s���1!�N�;�k׈J�+X��Y�����b�N��f�H�J��P&x���׶��'g��)�ml~�*ޅ�|�b	Eذm+��Ԗ�*��4
?�,��U�pp�åw�P@x��A� ��4��LXD��"�$XeUT���`���V���8�e�c�9�F[.��i;�v���x��:ᗃ�,�0��3�ߋ^<|����� %ty�C�ܵ���#V�j��#��Fn�?�K!����Ԇ?6s���W�V�~��'����1r��y����L!*V��ÿ3\��/K��w��ՠ���ө|�CW�c���˿Ku��#�Èo"կ���GWDKڲn��H/YxBg,�8��/�rٜ捤 A���#;���:���g��^�J�l阮��o)�֭�-0_-�);�>^&�m�3NZG��/; *a
Y�la�'��B�����M���c'�Z���!��E�W���؄5�O�J�v�=Mc�_���@a_�2�
���Dw��A笀'c��4� C�r[g��]���1�+����Q�)<a��	�$Y��ʡ5��������o|_��?�H~H�G<.��}�����6=�<`:~�E+ ɢݺ-{P��~�z.+�>e� r}�#��/Y�mX��%g�/�Sy_�9�e9�Q�P��j�C��\.;,��"֛OJ�ߘ�~�HLujl��1���3a-湿~U�E��=�vn_,$4�x�A�V�a���V�N3�th��/_�Jc�a�{��86�y���Sዐ�D^���3�5Hذ�9�['�(�0{'���C��#l��2��u�$%,󀜔I�K}+����EJ�g��G����f�UuV�R�c��d�%=��N�.�F���rY ��ޗd�R�Y$ǰ�Wh�S�|��x+����8	��N����Ht:���'�v]�49������l+��I�����t}��Q�,t��J���z�n&%��\������f�Eѱ�����q=	|	=����-�4@�8�t�Է�9!P�j鱑�%�>|2�_���ƅi	�J_����|_h0G�Ֆ�Bl8�$Y1�`K~k�2����8R��'�M��٠'	o�űC�Ĉ�r����W��^X�[�6�;��pq��~~r5��+� �k>�'�K��1q]J;�_ԍ�G��S�q�:�q��j�|m��/Ǒ�:{�D�h�޼Z��lzlt ��F�����$8�;gG���$~=��u�Z88��Ͼ!�/p�P��( ���B���^�E�G�+O	��[�H����ؔ� ���y�6�;�MG�pp{h3i��j�W��(*~OmӞ��@P��8���I��?K��S����s�k��\���|[�{��,��oU�V���b��e[I�.�Od�>��sǢY����)��ᅎ1x���H���Q�#�_���r��88�'��yUL�߱m	$�v����o�C%.��p�=#�5��I�6���H_��K�в�щB�|$ݗ��cѧl��u�\�쵋A�Yˑ$R��"�<,3;o�ł�_��"�o���`1��EIS'�SC�~d �5J�[�l0^��B�d��\�=K8�cyA�]ЖN����q���x<5�q$�|��yQ���� ��_a)3�Ԕ�b#�������� ��1�濲�	:YTmX�����W��T��{����m�-I縒����g��[r�ц������{cԝ��G����ہD�l���/7��_~�����B!j�q��I�׎��}���Ay�M�F�����oU���HT���v��6|I�%M&Bb)XR��z�}V��OUq�c�f���5�K��t��uy?�.;d$����yK27�Ĺv�Î´I�N����]��)�xj��%�o�4N;��%�J~��8|+4�s,���Mܣ�vN>k�	y>���B�ɀ�I���D�RU����Nt��.7�~"�T�,�j�Ou���d��s$,MN_uqO��NС��c�S�#أO˶E�{ex�%�-��2N<�������1լ�cx�>��qjD�7Rm]#[9�6�fzw��νmi�:���Ҷ?Q�+�i���H��9C}�Db�t�6����8a#�^�cǔ\���	��DͽF�j/�,�q멦��m����їm�4�?]��<��N�\0�!�>H�o����x�7
�C�BO���������L�2��v"��!a�M��&�$w����qIB`�6�y1%�Uc&-9��1���a��[wj��>d&����̩��$@Y�M�^w�그�����U�
�������3���W�A��	 qck��X��tJ싯{1��v+�)˞��X�{�Ur�8޲�ü�s����+5nn�$^���|(c�
����(;C�$�.��i��3�L
Q�W�R:b���C.Ǡ��'XJj���Cb��C�!��d�1S�������&r������?k�c�E.���;*�o�n�
J�gb������R��|S�c1��<"Q�Q�K�6 �*�Yh|�n�pƷ���؜*��I��?B�i#�E���јL@� �3���v��z� �������>e�V�z����Z�Nu#��_�M?�_OR7 %�G�Hn��ziX��������/�s*����������Od�C�EzL�̠��I��峛�z��;�}���j���^o�����?xPg�,z��IƙO�lo��O�.����N����L�+Xo�q�����<H"��a�z�K��vp�ńn+3�n�������g�<u�ڰ�tD磐|��{C�VC��eV�?�ڐ��v{9���C��ޔ����z=g������~�m�0�
�i��&�iڑ�Z2&�pௐ1�������k6��ey���+a�i�N�" d��z^��� ]>r�z�����rQ����X��U�nB7��|�y����~fH���|�ė��~n����^�ǁ�e�RO^��rn�tk�sk�j�P��IRB���%R�t���q����-��#�'����֗8e��F5����@U1�.WK��nQ\��DM2�/�j�n��=�����۝`o�"z����;bJX��!7k�.UDԊ$\����<ԓƛ�p�*/���-���l�='�$�:�M�f�k�;�1ɍ1��bQV���IQ6�����d�#J9�H8�0� ����ž��R�?>
�8C�󫀴��]�;�cj҈�h�����&�xaa���+�7 k�j[�N���|��p�U˘�ڧT&��S��]�0�����۵����=�YAtn�AN���K�Eej�gh"���Oe�]|�ۻ~�\��޽��
��n��?G��څftZ�D����Wf������	�:�8�(�Tna�c�}nM+�4?'N�������)0n?(^yghH�����/I
� ��Y�AT|����V�E旃ni�?V�ҍ@�͐�y��qGC˳wIH,PP}���c�P�>���l�f��]�6�����囹�z��^|	��JP�ñ�)������
h���_'���!6�{�։&)7a�䣽��R�;/�����`6w�Z���B���4���H� ܅B�[��� f��s�D�>��ڦ����,�.�݊��y���� �LXz��Kp�]XV&�-J�>}�[?�����TU���l�Sx����9+�8i�s�"xgB�J�x'z�e~a����ֲ���Tu,�Ϩe��\���ډ
���H��oO��f������@�1��o}�\_�h��L�w�.�m��Tr�FpF�6
����rU:`�k���	1"��;�!4J����\+���P�5N^7 C�wO�|P�Ngz�ߙ����'DI0(�\{&��/Z�᳜{ǹ�3zgN��w
pe2h� ����L<�y�7�ঔ
J����<���1���I���W��������܄�f�I��M���
�q�0��E>��q��YG���.�@E�C�7�oa'�.�o���Ǒ=�s�k���@�b�Q4��z}_�J������E�>��U���@#�i��yL����F���0'Q�����ql����E.�&����oC�p���P�ʄ �5?�)=�G��1Bs1�u�Vw�`$;wѯ}�kS/��,�e���*{�) �[�aŽ�<�ب=4<����Snnyhۺ��Cʕ!��Z�_�W���81A��X ���rJ���;����,��q~�џl`���r756}=�8�������z�!g�VK��ּ��;�f�T��=D��1��������p�Wѕ���y�2�q*_���FSM�դv�D��=6UK}6����7������YvR5����:E���RC�w".���Fs
��|n��Cܶ	�6�@��S�3���DQ��|;��|^K�%]��=rϿ2d(N@�Aj+�;x�C-(!��DoP��,�0w������'�EGD��f�9oT�\�snq�x�kM��F`&�F��t(�7�w�I������0!�LKKG���;o��nj���ǉS+	�����j�^�RsU���`B�2ML��`Bؤ��?���a^,�i˃F%"t
|�<����'��IΘ_)IV?L�,&�-֢KZ2��N�,��.��@A����>b�CVoR�}$��E�4�ꚟ��Z���p%F�a΅�m
�{e��x���mQQ���wa��#�j$�@a�I�i��9eH0vlƺ�!���A��n�X���`HC@���Gq�
,\����Td��:���U:��7�!t�WOH�c�������ZE�|Y{MU�eAɺ8�n�[u��R�Cʹ�Mq������O
��+�lK�f|����imd�N�3oE Q!� n��-��A�ٓ�����������6�-������]"E~�c8��os�(J���i8f_�u���N����A�%dl3����ʯ��$�5E�+��M�N��	B��!*.D87Gި�|j�(�5$)��,�!�W���ϏmuoA [e��
;��L;I6s(c��ѝ�n�(�Un��U"����|���������a ,?�F���F.E���*�?_��R���M����o-@��1�o����������hc���#])D�r[��wt�;e�87W��Ξr���P�w��SA�3~]�`X���M�й_�7��W�Gq�rG���d0���� �a q�a�ۯcE#�M΂�2�O�]%�Hƚ���ށH=7�%8�Lp��ޝF�.��!x���!���^kw��(XB牬u�̀S�1���u����DG+&
�
���tB4� ��UH�y3���T��V\�b����XN���^�sD�;H��7��QXA7��`=��I@

�z���n�Ӫ�_&�a��e6j�7d�3�:h�3j�nvr���d�Q�L��S��J�����e���%����ڲ/�a��
����i���~���YS�ɬ����7`yR�?�b9�A�ǿ_{�>���F�'�+I��� ν��[O3�2��:�4Vi+t=d6ch�	$�/6O2(a�Ï�,Ջ�N�E����
x�bv��B%�J�!�SX)c4�����MK[n�gB�#����y9�ܸz*p��^��,�h�F��~c{$�Ɇ���?�EF�����/���Gw5��Ռ��v֟��+�FQ��6I�`Yc�Qgj�6q�z�toCXm���-R%�0z&��f*H����	 mz�2\~V��$�-P�!˧J8䏙Y���!���km���W�T�#�H���/�� �cd��/x���9�$�vxb�H�N�?I���/��$�^��Z�M�Ϝ�t��x�h�΄�J��w^]�ĳ^G�d
Os��N{�H���ס�i�=BJ(^
��xf��~;i��r�ߧ���2����]�$��C�=k2S^L`�'�2�դ��t�`�y�	6_�k=OC���h��BJ��@�G�I~�%���3޶�aנQ�S�����n��2�K��T���������F�!%�E�间&�,	�dsd��hEh"���]�qZS��/�M�]�T����V%�EA����E����_S�-KH��0=&��d�dC�H��"�%�N]���`\����YG���U1�6�;�T cr	��5���I��7oGbu�3}�#��;��WT?w�^���tI���UG�Ɛ�%��-�}�_+)�fj���O�-j��(�iF��5B�~9�}ݻ;�C����our�G�� ��fbgTQ@�'�=1ߠў��gT-����w�3�2H�N�z�Y4���b�o)'(��L<t��N��q�mh w��z�共3A��������5��p�RԚ�y)J2�o��F�>7tdAk�ݙ�0���S�J��oz)x",�.����-�"���f���լS�&����`�H��¢���M����j&��OG����(E�z�=����3�A���˺C�Z����6S�.Vt�#���/����))&�����r��ު~�L><�`��8�[�ƞ�-ϓN_Y����qOF*/��&�E�T�;�S��
��j�Ϸ�Ds{(oI�[���IU4�~�F���(l�Tu�gB�m kn�M�,P���F���U�xn%Az�}F���XV�����K�˯��`�0֥����u)Ѯ�#������:�n
���_��S�?��7��NA�O\8����nw}�q��̅ȋ"�i`�L��s�
tD���9���$�*�9'X��p��6���[�T񘟻-M��5��i���3�E-f���
==���ʖ��	 0��:�{�!�֥A�`��:<�|:2����! ~����,i�5�9]<_�̇	�@c9D����������Sø��^����&��fD�B�P?��[�����L�~ؕ�J+i	�IN�9/���j�ʵ�'��^Q>�޴��\��Q�����0i��,]'��1;�'�՟V-��8J,E<��S+�P�T��G�ِB,���z���S���i��I�db���<��"/�Ka���ګi���v�F3���)������.���Ż��~4�6���\u`�#�#�wTP�<�D��7(""��D���xzf��q�Mx�`q��N
���@1�J(+`�^,Z�b��i�n�5$7��r����=w X�a�0@��7��� ��Js�R*A�
��<����o���O7��3P��w��8��]�3�;7���i�����I�RcE�`��3P,FO
�(5UB�*��feӝ8���Ehc�w���j����JW���R�b۷��-��*Y]�S���+��.G�pn��WU����)�`|���EcH>^��I#�����>
V�_X@�fN��)"����~��q'�ZU���}�s)���[���}��*�?�+�]+����>���w��4%l�6�?�������ݜ3�]�~��LM�.W��*���ViPSKZ)j��(|����09L5����������Jo��Cm�+|r�̰3J8<�:���,;��M�̏1�*9���n9���M�]��3�ީy��䑅1[�OV-��:r�m7�gS~�xך����J�Y6e�C;d�?ywh�����$B��|1��&Ț����!�K�غ���f�e=��'�����r�X%q���~�{�i������ �U�=
�`���g����S��l�(1;L��N�y^"Yv���QT�:c��;��r��p߽�1|��_�dzL��t"��d7�r�x��i�԰M��v�1W�p�q�X���	J�J�_�RO�H��Zx8���6��f��}&��Y26T%�aK��	��{o�n�.�+�8&4���w�$g'��&���N�:-I�y���B��Ԡ!z��c���ц�ә|�ըf�V[M�y;��	��vk�a(�zC����9��3�]�2Q���dY�>YO��*�&J��ކ%�x�_-p���E��d̽���W�����N��{�wmO�mgF���m���{��]4��Bz$0�c�)<_��a�A4^�I=�bʧ女���/�] ��Q��ߘC��Ճ�qa �?�+����j���Л�p�4�'����_�������5;�J��<��OIeU(Ȱ�1�:k�t
;M���<�A�t�@@M�zS,��([5�ֵ(5-���ԡ�]���(_g���5e�LYٸ_׬[��)������[��(��<w�b�9W�0��1S���x�v��G���m�Z�d�����8ͣ�d\���j@h�xF�q�d#h�rJ�ݓ�{ġ��"j�]�dn��#NOӠ��x/�c��Z�f���Ta��GϜ����<�7`���Ѿ�@I��k"5y��X3GIŴ��T1��s��s���Z���2k9!��j�i3��u�5���������UB0�i�m|�rA�QEj��>=��=$h���hJ�Am���/s���CϞ��(B ��n{�IW�}6&BC�&3�8�TV[̡�W[�T"�PG
���Y.� L -I�yFO�!�¯�l�L��9L���%=0[s�d�)ѫ�E!��ۃC�����-�`>?��k� f_��V��~Л���9�Q�P���fb3��z�)��w�ǚZ��.�����vg~E�AV?1����B���κ��D�%���(�z=�wu��L���Wn-��օ�e��<ӡ��7�4��f�R���"���0RC���<�SI�/g�|�Uk���+�v�w�����
�Q�4F-/̌�0��U�ڜ����4F��J�@����l�lm	ƿ�mdCS.�LT˵`f9<�\���uq��9D���0NG2�L�����KYq}|��5~OA�7qq�Ё�T׊@����烀�����	Q��Y%4w}Q���D�(�Hjۣ��dF�RdT=�-��R"��Vg��z�ǩd��&Eb!��7�K�T����_d�6+s� ���P}���E��k�6I�����HH/�j��,����Uy>W1�L���'7w�s�������h> ���,,XA��^�����f�`�P^��Rw�Mr!]P���W5��M���o�/�~�*v�d%.4����Y��|�Oo"P��#�b��DX~���#����(�~A�����&�.Gu)��M�'	��]��+��:,8�䔿�1ފ��V	gZ���`)�K�u�ZԸ�g�)+�����N䝻���D�j����'|�/��^'�1x����J��6�b <b/�\A9�\N�{�H�0��F4CZ+�|eJתFӼODZ��=�˶[+��-�Ê�&;or=r��e�#�$�Kf'��;���ȍ	O���NO���F�p�P�+��"�0S�w�z=t��7Sn�-���~��-�[F�W�^���
�.�尯�U��VM玬�×ڱk?7gJGȆ=���ŗ*Av��<���Q�L%'� Y�p �1��V@_#�"M�v�m�e"+�W~�)���ݭe<�'��.�B���F��Z~�k�Mn�/&cur�	�>4NUc$�-!��;�ݯel�Dx?��c=#��Q�^Ҏ��-��!brIֻ:C�˸HُpKFu[��5�bH�0�X�%?�AH!�ϳBr��Б����f�a��SI��C	%7Nn½���(N���cT{�rr!v�UҒ*Oo�����6	��uQ��[�k
_7���L���jdٵ�w��4�l���?7-	���^Q�67����	����ר��m2�S��LR�Rk-N�܊%�t��|(�܃D�y�T�-���\�PO
 ���q�Vr�ğԖk�S@��*lF?)g
�Y��A�yX)��𡆐�:�F�Q_J|60N�һ!����o(�ѣ��Q?~�B��� �n����:ꉱQy���c�A t�W��UM<��O��(.�O��IK����Q2����K�������[Q�T��������d���IDK��T���Ǉ���p3�b��=WaqO��ɮ��zR-oh$9�D'/�R�X��-�p�W1Hx��{��Rl�{��l� 9�����<��&��RM@"��9��5*���Yx|N�Z�t������/��J3�ԇ�(.T��S����/>��ŏ _Asc�A���O	� }�����j
��I柗�:�{,!"��	r��?�Ii��Y/��ٵ]�:g�_�zյ���l�@ff-?������UM��(AH�4�i� �>-("B�YWq��9ܬ:���CËK��;�P��]J����n���ͧہ���y�ú����P�
[�tm����ڒ����M�sT���Rb����1�A��u.��1�)x<7R���g�=���;0db�%�s���m�o1Cz�_|_����t�^��c�Z��{�ր(t��2��f�yѸЉ�;����U���@�;�P4����v�~
dx�Q����ڞN#�?&�d��Qd����=�hA�k��\Ci��#@��ݷ3@R��#Z�2s�Z�E��bڛ'�|Q����u_!�-�L�[v�;�Y�O$��V5,�)٬���%J��ڰ�^"Ԡ0��@����9=����@P���2Kq��H&]y�e&,�	t;d����<,��������5���[ʆV���%���f��~�����,0X�p��t�1��?��~��A�I��CV� ���xP4��k�X�nJ9��U�p�����L�?��=8����J���,�f5��GWk ��Ϟ2BaE�F�����{U.5����� ȱ�����e���7�Tǟ$�ݥ�)E*Er'ya�|�"T8��|0�c��Sjc����,��K��m���#%m!X=�����Ȑ��mo���	O  c�X��k���������f���]����c���K��%M�g5�]Æ��_j�z\�mp�8΃� 1�)T;l�~9՘�-1������ #b{���r����?E�	�ol#�+ar9 �'��N���1\���(�{�G�����Kf����A�
�{\#��|��*$~�զ"��v8KiP�ֵ$���ă*����� 5ckz����D�(�& �D&��{��"�P�G�f&q�/���ui ��(t���N�6�`iH�7�\vWw�	7̩�l2ޖ��[��:�Hc��(�>/����G�	= ��䃷PRL��AԿ 8+�U4�^/;����#��K�oT�`�I�̆���C�#8���o��l=�0L3��U��X�� �A���,�{cZ'�$0�G	-���u��LI�Ǩҿl�G�Y�m�{�aF�-�����kf�vm��ƾ���>`[��[�f[�VUe��o��8�N��_3�	�t��yA������mxT��$/�@0�V��+��=��ʟU9j��Xa}߀u_���o��2��c�E̞8���n�3�5=fגZy�1��n� �1BYRm�)_[��y˦[!@-�%�l�'@�ea6�*|�`\��Q��qO��2��+��� 	�Ѷ4N/�b\c�LQ��W�Esh�ʞ��bݐ��kL	۝�'��Q��G6�k<�Ҩ���h��[���
$�ɸcmc"�u�
+^"�.pw�%1�;��&M;����MK��#T�f�h�K=Ni\��櫽��q��a���G�<�U��Q��e2	�[cJ8�Ӟ~=l��k�v0�F���.oS)u�z��k�~i\�k�jB��R��o�Jpq��KG����>�V�?;|��`Z�P-*��*�ĨK$Y�p~eŹ�R�g�M�#����;��BSmy���O���<�oiϊL^�����x'{�P�.��N�z����`� ȱ�,%��`��ʔ������ଶ��l+�D׸ǩ�,,���^�̀��=��y��g����+7x�F�a��|�����̾R��]pB[����%�3�#<�|���=��w/[ƺ���d��3>�*�j�|�O4;��+ ��Y$D�;nG[W42-�F��,u���/���E�JbY��2��_fۤ�H��e��2$ ���B��Q�ۚ?���U��w���c~aGĻ63ں&�'�<;���G�	�����hضM�S9�S#~�u�����?6�ná����64���!_{�{�����a-O�1�c?c�f�낚�Tbn�c�Y�U��q1VZq�l���u��[X�/�z׹�(��	�Ȣ���O:j��?m��h~�]��8H�Fg�K�j��x����g�~M�ܜ�Kr�6?6�jAXD�����T?ugA��|�/nxZ�g*�L�ۜچ�i2u�>�vΜ�l-=31�~�fE��q�@/�ɳ��D�d��-��߹�s�$2��*����m�)��p}	8����Ǧ7iD�g� �h��eMYk���kPu_y��]?�t#u-�C����j�:�������įw�5�Y�R��cX��I��l�n���u\�=���v�dw�I�a ���)S9\h�l��3����)�P����B�%זF	��3C+��#��j�����"5��Lt��l�M�Bw���@����� x'�t�PK\;���J��"BL�Q�P<��yh�U�%}�RD�8�� �V@�H��������R�Q����ߌ���q���1��^j�g�Q6�Aa}_�~��T{�����:������{��B�����v3��ip~����A��Ju/�w�5�˂�sH�ֳmdAw���ڍ�w��7P�������<��v��RD��O��!�x�80O�?FC���z��ȤH�I�z�q��e*r~���:m���GU1�u&����Lz����h�ԴgVҗ���(�c��w!��J��ߞ�cl�zX��J����CWr�'���?�)=z�H<���595Yx�w�tqf*϶;	��Y�����l�3U�Iv�D2�n\�Ň�r�Z���v{ʕu]½'��[��8HX�YD��X���B�� xԹ��sL��D������y�Aw�õ� F.����'*�u�sL�	5�c���"��/�J�;��;����$�4������+a�dQ��[�A�de.�Q�뀣�]J~e0uǡT.���ϣ �r��ב�����TT��s�0�D�ҿ����C֜4��ծq���%hV�Z����u~�C��~1�ԀS�,4��	�!����\my�/䧽)l�I7��tuB���R���rR�+i��@�(�G.N�#?X�����2T�]8�.�Cb!/x�I_J������dQWZw)�䤷a7/�U�I�
�"�7t��a�h~�UQ�p�F��,U� qel�ؒ��u�$��vH}w1:�@s��p��E~����>C�[Aє�	m�kD~��K&�9(RJ�F{��T+�g��Y�#ex�\�R#���e����\�(�&��Sl�	s���;�Q�Al�@Ru��zeV�����O��	|4��z�s��'
x2Y[���@��VxYq7�P�#��Ow��W��i�c���P�����2!��.���_�D��(B�`iF먚]{�GB^NN�R-�SU@p�ƛ��y��Q�B��}fGS��F�s���f�b��X	0�<�ҙ]����sI����IF�K�
�_�eDd_�OM<[�w�O�*%������_4���\Η$Sj�3���G�Q���D}�3�����BG�O~5��91M)�>b�o_�<�-$�nϘ��j�u�c!���4Aq�9���;l����q��3����>�m��_Ĭ�=�эD<����qH]��<�;��Z}��,Ms����d�?���\\6ӽ׊Ǽ����X_2��4>Qٖ���z
���hpoօ��ע>�#�W�Q����93��ֹ�R9$\jm%%���Yg|�e�J�.�%�a���#�y�/��-�$�i#�K�L=���b��D��Ӿ�������27�up�#�����)v��i�����WjT�W�r`oEt:��&|�I���7af�<�7ɜ6%Ȋ���0���q���*|6��5����t�ċ�:$ɧ7\@��W�䮹����x��N^V������-Ɉ�Zb��u�{�-Yv�a�ަ���!�P�v8�\'��ZwD�������-P{$�9R7�K�Z�$�������	�8��27��+����0�𶌅^�&Ql�K����;�������X�+�$���#Ϧa�gt7��*h�����z�,��}�_�-=~�
\F��z��rƅ�dܢy (no�)�ɡ\y��3�E��de������x񅊎�zⷉvɀF����u;v�ی�^�{e�Uڒ�<�Z����D�N~df
j�L�Z�Cc��
iU	�F���B�%��-�E�����~�t/������I�.���gj���^ec4��88�>�Wdx0�ZC��W��$��#&\�􁿕z��MZ�a�C����HUg��ȓ�L�igz�͆�{���Ou�&�'I ��Z���K�l��Ⱓ�ǌ{�ٱ�⿅��4)l�|���,��O#�r���R!䔈\�z��QCb=��@���V66_~ӝ<�Pi�G��٩��0�۝4��g6�}��|�W�y_;^�0��S�b0�^.���q�����D�t��5D�'d����i�׵ꑛwФ�u���z����H�g�����F�T�(��D&/���P�&�Ӂ�����)#L��o�@�[��{��n���h�t��\=&���g��3�G�Jq_;��[�%�`���ޔ�hD��eN@6�#�� 6��O��+ZT���ӦA󋓬LM�!�UN�`j���3�VGAd��n0l�ʈW��R�w[u�5���-Ԏ�TA�T�N$.j��4�\�Ϗ�A��e	�!�-�pD D�,��M}�-&R���Ц������f�E�K�P�i��
�l�sE�f.Z�)4�Ǭ����K�A�MP޲�78I�i>v���F�YVy'��'i�
�����F�`F�tX/�Ë�h(
&��r�WO�6Ẕ�6��4#:NpM��AY9z���ML���>	d���jqHJs�����E��-u��Eq�y7�����_=��g.9i�y�(<�YW}�R�$�i�nv��#���.�NY���̴�D��H�C;��A��8#�ܐ�*�Ǩ=�	 |�2���h�D:�xP*H�����k�6�w�����6�*(�_ST���N��|�}��~C6>s��o a��H�����t/��{6��A��N|o�w��n^� `�I(�K��~36$*)퉘�������y�%3��=0�@����<w��Z�\��@p�ь��<��1� �,B������/L�<��Wr󳺌F3"�����2Ǔ���Q�8�W�O݉gɷӘ\��&�H����K'�6u�&����`�-���M��J%��0;6(_�f�H:������;j�$Ӏtl2���u;1X�)��s��QP"�GPD����+����H��lm0W�t�H�݈R:Af/ru�=ҹ=Mzg�N�[N�R	��{Ϸ�Hl����㛟=��b�cE�f%����~�ل���\i�l��P� �0D��v_��,�$XL�2��e1i�J��sDf'�n7Y~�*�f�ʶ�;Ȱ��-�,�p�<;%,t>�M�r:�=�[��`���8�A�������NQ��p�c_ZM�I��r�<���{9�[�;�-�+tn8ҍ��\�+�Sw�=�6��a�-{�^$k��?e��iaLXb��ot�=\���YF�:��S�h�c��6E��k��ð�8ۀh���^�Dh��v�;G�[�8*#5��{@�{o�ۺ(>�UgKߟ�)#ȂD��������-`&��}���S!Vu��F��7IY|O�c�C�q��.�
ygOv>E�K�9�N<��{������N�@�pe��r�;��/Bs޾��`Bs�x��k���W�p�i�����3��X���)K,�uM�u:�A�&�@j�-*�ר��"S�k���PB|��)����n��:�nն����U�f>��7kv6��x�_鲼g����"8��m@���T� �0�-B���kE� E`�P�1/����!V{ø�u���W,Û�����9�w׿�-���L+�,R%��[7����@!�tj����HE�L��T���n�<�@���A-������C�𴐉OpkWpp�65�S�zS(ݳ�˫���+�UQސԠ�'��%)(��H��#����:�e���r��hx?I@<�FS��L���	�񁢪�/��Ú�I�Z���T��Gj���y��wi:��鍻x����S�r���>bN���^F��~�%d�މ�x?�(y?d4F��@O�����Ry�D|�{|�s�qKهU�-_��L;���vE�'��dC���v\���>	�4��QY��WA�-�E�5�e�΃���}���xY��.I�jP$����G�D�*i���D�^�Ѝs��$ͻf*6�K*#�6���Q�?^�t8a��W �&�ژΌqi\��/i��p�>N�B=*Y�^���ʦQ`���R�霹��"�c� 
�'�W�)�t.�d�tȞ-X/�	߻'��q��9�2�iQz�\$����y5c�s��-�ц��y�C����r{|'�pFz�\�B���o�Z��|�iń�演�)Pa,^8G:������L�K�A�Z>xw<��[�oF�b��&@E�J4�-ȉb��_��<�k6�B�ㅐ.5
,��有��+�D*ě�p_f\�H#O����e�-L�v�y��!r7-�!߶�#ۨ(�.#���W���t��]�����n��h���X�Ū,>��F�t�]��ݎ͵^ؒa5i��L�R]!�]F�ۑ��e��z��N�[S�b���d��+(�"��1�����M��*/�i��g�jtUխ�f}�]|=lQ��:j~8�HV�E��6U�֊�Q���_Qoe�����yѳ
�b��5�'��	��-wF���Y_��WCJ��7�����6������#��""���vMyC�����k����!�=$Hb���i����`��_-��|�n��h�i�Ivr��z.@6�~=f�c��N�����xG*V���	l޲.�tT\�؞|��!d��|�ǠVT�)��̳�N�����(^~!>�b�HB��}�ǇQ��r����k��h�?��>!N5�W����}�7�i���K�	u(�e�����k�П�E"+M����2�a�������SB��(S� ����3�c�#���y�=�ojUH,�3�����f����3�-���J�v�L���	�X��ɺˈL,k8t��;x���/�����+3�ԗ?`)�0�: �<o�BL
�a.�n��(��]�q��FG�"�<�(V�~�&1�88�4���l����Y8�A�����zs�~�3c%�3�L6�7��y������=��{��6_�|��i_L>җ��7���{�r*�S�chZ�Ə�r~a92)�᧦uWF��!��g �ߨ��fu_�n��7��oAd��1�1ޟժV��Rd$�>.u�Y1�5rX-�&�޻�
Y0B��n��	,��w�*P����9�BmPC�+�K���?I�9J�-�,3��?j�ԓC��Ƈ��X郖 '_��UĞې��S@�����_����w��,���hY5�3�i�Hɿ��	u%���]k=�����.��*%|�D�����2�$�f:��@Y�8�"�3���'>�X���p�9�k���a1�J�!��G������`��ƛ�'��S��B���Ѡ���k:�1��ã`��IE�8C����=$�u�R������s ��0Kӄ5wj,"��bɢ¶9 �Η����X
�2��|����%{ ��ǳ��%����<EWӌ�,���u>�M�F�k��E�9,�jd,��XMd�3����^������&�\eX#����'�祦WD�� 	gQ�YB$+muY�����������<�%�4��6�	(�z�@���Ӵ����ed՚.8�sˈ��"��~QR�_�=�>����/\C�
W��"4c��)��n��ڝ,6Iѫ2�� O�S��{�ѱ;�Z��9��ʤP�W-3���Ͳ�����v�/���_R�$��T�@	*��i���䧐��H��N��ju��$�o��ԑn�[�=@�0uՉ�3�j�׸\׻���w��1���|[k�&��⻽ FӀ��T�]���s�4f�2*��X�[N��F��qu0K���c�;���@wScÛ���&�l2|� ?��r�h-u�߾M��>D�F�IN��5ѐϹ�s��p�UnV$$M3}]���ݭ���Uq�E�4\���[���^� �v�{�E�<d4C~���Ȳ�3���J��|$��#�Y܍�7����
��0�1[9)
e/S3hBY���D<��h�����Ȟ�����8i� �M<����3���K��\�&�}���A��Lb��?�C͛b��5X���3;<�.��#"u��ɽk�n�}O;�o�0,x� �[���`��6-��
-��6b�7-z���c�HVj��N���%���9����R�`黭I2�Lu�5���H�t�b!���a�A�Jy��fَ>9*F �jd�\�s�ƛ�k��>{J�v�&hC��՘�^�)L/���17�K�����^�g���y���4r�AGCs.�A��a�S��|���}Ҏ�����_h��Y�ի��1ZXv*$}��=Uh�TR���TcF���i�mq	w�U��Rm O�_�:�.b�~����u�1ޠqJ�j�2�@� X"�XV<������QY
���Xɓ)��~c���獳��؎���8+�D�$%G��KZ�uK��|x�p��)(h�6,Z4�o`!;�oCТ���l9淘2�);D�l�F�T��d��3��%��p�\^\�VE�"s7�����1�p̉�����VG"��ho��ٰ���Ekl	>&XLX������¢m��*��q���l+%�+K��u�M�{s���: ��e�H��]�3O��'Ui��u���L
����j}��ثX�gή������S���@���Ĩ��WѠ����:c�^Ԩx�T�����=��͗��V�Ƽr��{�.��@�P���[�HU���t�R�^��r��]��ǩ3��B� U���ô�CV�S�H��sy��ɳr�%�e�f\�@��L�@�}�hI'033,m��Oi�ȍ���h�L�F��Y���o��+���&��� ������{!9�Tk�+�Ќl���O�"�K��n=RLlqKi�W��z��U�<�	6fW�n1�8t�g�,�J�ϱ�1���e@���Z��~�d��8��.�"1>߮H�
�)J��w3����"j*��Y�?����
��p��1������8�2��\蘏}U��I(��yZB$��C|��`i6�B�a#y��GJ�O.���.��a�#��uMX�)�is�+�wb���͙M���9���|Đn��V��?X���2}�a74ƷnO��)Ef�B�Y.]����..8�g�V�^a����"�u�	�M��E�pɉ���2*��wt�լ�7K/��98%��s�1u�J��ʏ��;\	pں��S���6�h����
ܯ�&�#���U{�1�{�}R����1��� ��8
z��Pk�I�`i:��"�qN�Ħ<�5���.�.�x���-�Z9�G�OU5	�DM���H�9u�U~=�L����s������u��hцyr��t�7l�O&��o�nm��>�zQ+�I��c�Q�v�O��Ċ-�Ӂ���x�lhBU�Ev��߮���^ 
O����؂������ɼ͘A��5ph4��]~~�x޲bO�8��Μ�Q�i�|��3
c�>7��x�_����۔�!�A�Q����IW(����݉�A�M�U]�a ��IH�o˭
qv�V-������Ks�f}°�&�s6���({��X6;�=�:J�(�c�ҝ�lc�/6�g�R����)�gT�[B����vr��������R����x�#��w�Ne�ۦ�4q+Rp�C<�e�t c�U�ܣ0c5K��F�W�|����s��ʒ*���Au���y� ���H"�ew�l;�,�;I�0�h������_�kZ>F��k9�g�4|/�Ot|��R����v��q(P�#�l8ӽ�l��Ѥ�����*��v�{г2��x�'r���G�#�0jLQ����H4��U5�=_�����J˔3�$ �+LB���9���K?�Nj�蹀	!i��DI�C�T=V�g�S�<Q��2�,>\\k�'�m�,�j�9���bb��� r�P�UĊnsqA�����d�ˁ���>(��;�;k��Eμ��D=�Y�\��V�}�&�%���������?|���w�X݅_��t$�-XϜZ��>:��Bo/�#֮RA�~�+(m��Sug�Y6-��h-���}}�y�{r�!V&�Oئlx}l���r �Z���C�O���r�ï��Ƥ�j7��8��I|����N���r4�|-�{}x�f�B�q;��xz�Hw� ��|��R*��t�y%������l@[|M n�
�p��*E���;Ϟ#$�'���f�q]��6ׄ��9 ���6�ۍ�x��6�xQ�d|��*Q�зɭ0�*}EEi���i���+t�&c;9)DC�?��mA�)�l���~����U�J֥Z~
�2�������̔5X'QN�1�����'�vŠ���-�r��6)�^�%W�/��,Tn����B~ ��,���rӮ�`�"Y6���rK�:GN�� jˑ_{v���kNE����@�NGV���E����6��frTq�`��H��2�H�gC��>� 20�[��ix��'���	saVZ�:����X�[ЩG��Z�/<"���u�G��{}�.�|�bKگ�����xVD���A�:p���<��L�!'\�Ūs,�L"�I�U�W-W�!�]K�)?�"�`�?�m��΂T;E�v��ݰ�2j��:��,���N�ӣ<��8u�5P��`]Q����wO�(���ؘ^�-t+/�j��c�݂W,8l�"�D�����U��8Kp����Uɀ�����y���
ձ�<�U�|}ᕄ��ޠ'+�n�LX���\�d5����d/����b�
�?��ckĔJq���=�H���Z���vb>\�1\���=��h�⤛|e�G6�>�t<�#�&��Z�N7���Z�^��,JFѝ����F\�eEh����s�q� b�U��j�f��/�:d�LyֶH1mlB����gn�[K�tS�L�+����v�V�]%�~�Kv�[��D/x�<��K(��(E��ܶ�^��ģ'k�ZUn:T��fO�iv�"�vR�ߩ�H�����l ��T��R-���K��!$4-$/��dP�$���C{x�D���"�T_�X��������;r��9���_�I��Ω���|�x�ٸ�k��s�P��19�t@�J�k�Z��<��h��W���r�C�@�}�ʚg����3�?!\%�L�ji��k-D�_p:ܹn-�h���ʾdE�@.~���n�
"��蝑����抱��K������AmdW�'T:�#���<>�ތ�$ȣp��+I��F�gwg�l��2�{^$�1��6�����3��y yڤR�� �iY�Zf�z��X�+�>I��h�pim{B�N2 ��a����rhj�]�pev�L=u�sSk[X� SS��X�J
�1�a/wA�u�\����Ty�˵�i��2���\q�-�K-� X��� ����:�=X�i�)�E@�X�:�[�qq!4�MU��!�Я�~�j϶���+��{��mN�Jg���j��kmMiD��|AcuIޫ�Z�����Z���^�%�;m�8K�9��|)2e�&�'ÁUy�P��}żS�A��#���oQ��#$ ���ۣ�Q���E�',7��]ԋS��[k��ɪ"��u7�w��BXH�?ɭ�#4��c .wYt��}�*N� �r9���];���8Ә	[F��0���a���B��_����0�F��p��y�8c�n��!�Fd�k��<l8����At�N�4���g㵋���_	�(v�Q2����o�{�C[�t'��UPoVc�-�gX����"�߭2c�:x�[�v�4�����s�?
�Os:jH�*��9@Mf&?�y��[]{8(�KMJ�N�|�� )��}���-��������
�F��*x�QH;q�aI�/;n�Q���F(�Vh73����"뵎�y�U�kly};ȸ��I�H��Q��K�����*��/;{����r_FS��H��V뇠頌�h�&bh�����e?�%��,Z�C��,g*��!�A�xG��*Z��w�B�ܼ�r��j�=çݲ�s�a��͏��Jn�4��²=�P�7��>��*�l���{��i�q|�f6\Ȱ٬�+%v��R���������l���|M�f�
~9�o��^���x΋u�c*'�:]5�v[�i�]�t� >i�=���[��kv��%�4��3,B�_Lmc�|��n��h����@;R'e������e���Cp߭��"��
W���]X��d�j�X_>$@����ԑ2�`�Fʗ��@8׀�2��;U�Y!�_��uF8�x@_<L�G���(����<��ŕ}Q@�Z�QD4+,�7��;����~^��[�u��Mͪ�f����啻��6_�Pd��3����yD��
�n���u�;Jc��S*�mA?$�c:�vfU+퓿� �:3(ֳ�4�0�R�@?|=��2������z@�����t�}^���H)*s�yU�ߢ@�pU�e ���/���D��d��7.6�OC�\��O0^,Fs*���Ɲ=݆ӧ'�l����X
Z����U��co�3l��:����^N{$�7�;����v: �r�<�*�$l����3��G�x�VK�T�BU�y�،ܫ���]mTk5!��:�}��e*�J�k�Aa +���,����.�n5l�
����c�"t+��(��D�pϛ�&EN(�t#9�fy*%��]�=�^�
�oe���"��k湲�4�Jݽ�7K#�c��xZ���"G죵���S�;*����2MX4��?>5�wa��
P-|/3��Nŭ��M��q��vo��b���]��LY�B �ҞB�H�X+}��U��/JARe1Rm&�ć�~�S5N�&V�+���Ď�����&��U�;\J.�ƼgH�Z*5��P1��2<��>U�-Z��%W@D�w�ӵMu��,Pz��I�T���f��Ѱ�xe�l8�*u���u�����*]o@�2Ӕ'��{��@h�)i'�A��t���\�<�t0��[�'&�h��������{�z6B �O�"�}��r�o���nh��\�]�z�z|��!��t/��dA.�<����f�SǼc��pZ��?���(>����Z����QE��qT��T]��T���m��OT����\k/���˒������e����.e��Q�>q��<��� ��(�m��e��m���t�3S[3��i�
�3� �t�5�\l�?���l��4"��������J���Z*<o\�7��K�s(�t��}�[�<~�<�-�:]�2��f��:#�ٓ0D@�}���y��I�(|.�+�<�f`d2y"�����׏�������ɫ͚g���W����9q���|є�+�;�j�A�6o���zi�n|6&���m|�T{��}\���O C���?-�1����C�ϻ�L��̨t*a��
��I�?�Ht��"(���������j饏B�xz.7�͗�,G�>�1�QͲ-/�PK}T��Y������10�uQ��H1���$��׆ *I:�騭�}���k�U
����rT�>
v��GC��O����W�aTUꉣp�c�t��~2aG5 �� �$L>S��O�zaA��z�0�*DL�e�ީ3ǡr��.I��ث��F��Xn�S�_��x��#���[%6=�g�14��F��*^V?9���/��O�>�L6|R�)/��_R}5_�-u��L��ٌ+׊[Ʀ�<@'r���˚��$tn�$�����!o�YK�؟7P�.�cI!� �!)�W�Y����N0��<��O���F�-E��, ��j&�XZ��j*��,�*R�1}ܤ���,u�aZ�0�j�^����NC	�_lo�q�LZ�%i�GN�u�F-}M��0F�X �d�=��g�5�F�K��d\
}88B�|^����a��]�M�f��7���|D٫ss�tݗH/�h�ۭ��{bJ̆��¥�mng�x��+�[k�+��Z�ՇREc���׊v�o� ĕ�>�0��(M�݀/z}/G2�@�)X�ە��(}f�Kw���d�){4q��!����K�/t�p��	B�v�FLh��r\1~�<84{��A��9�\��5�K.�=�fF�oP X>j��	))�k����(��~����{/KT^ۤ���B�ְs/�T�n�n��󰁍`۔w����ʴ$e��;	�Pʼ�$�M��X3��W���q�LR��
�� ى�K=�	売?�*W,I]�\�[�m� }2�PD�~�ߺx��!�V{�������D�8�]�k�)� K�����U�D��ł�hM#z��CPӜ��c6Ӂ�?�%��2f7��ۙ����4S�(�Y���}�����@X��zv�yջ�0k�lm�1�<fn���|�]Ss�Xs�Ԡ!����hN)��bj��7��.�Lq��s�N(�܊��0�p���4���.q�{&eJ�8�`�7��`��2�y�9܂����t�W�~���!G�Ԭ���b7Pք�8�s�G�*��^_�U�_�8u�
Yn�mq�0�q��v��:��7��D����dް��j��xm@�rB��>W�!��r��?��5�u��l��S.�+�/Ѝ�Q�:���������Q���R�;�MQ�^3��]J3�!��c�7�������o�̉�E�W�
��K����ن6���3#B-~����d���Q���ج�xR�S�u(`��Ġ�|(*��/"�O���~�ϬE}�%�5�Y�_��y�<����z=��=���V���h�x���Ym2�p�:!�\�Ȫ}��͵B( f�i�Xd����V��{�\������fO�;���4?�
I-�8�����b_R:dӋV�h�bw���&x�N�!��p�1)��E��]�}���m()�H`���(�	�u��;aM�C��D�Cf�f� �t;�p`�%��L��1��� �W��>U�V�9hiQ8�:H�u�؝�z�q�\X�0�5�g��O���)��>�q8c >O��tD�Q�3�X3�t&��+?v�^K(9g
��7@M��a���_mL@�n���F�E4t�[�uJCG��!Iߪ��`)7��,iА�鱼��p�y����EO���:{Z�t)��Y,'F8ɬ���x4 ���`i�J�~Z���Ϧ�29U��_@��K�ۼmٽ�~�$�TY������J�0^�L>K�����*!��Q<)n�
)5q��VK����.
��K�.�4d�U�~�"R���ܙ�=hÃ=�#VF,�iuĒ��ߘ)Z��YB��	M���Pْ���f0�@�R����d�J�]Sк���r�i��>I4ay��=a[�?��&&(q��ۢ8�=q���VyC����o������*�'�R:��;�b6�.��`�����"d�g�i��b=J;;)���5|ZY��\
��i�"����0���~חS'#�n{p�f���Յ�B-G����)�Ѓ��J6�m`l��y����0�m��/u���t3x�k�����#$~C��Q�Zv�GA�Y��(-��~�3g*���
�x=&��:����BR�u{�K�f���զB�lǊ7�6-�7���|�fk�k���v�x�h�ue��]���@	m�&�u��5�(�� �!e����|�p��#�b��y�4��L,p�0�S��[���F�ޖ<0��ﴻg��6*�F��o3��Z`���'�)��_~�ӂ E*re3h����,���^.���ly�������k��$ܞkJ�o�~Y����N���F8�cb�Bg��{+<W>?�rX#^�0��Ĳ��3-����6�|�qw���L�0ľ���zZ1�*�7.�ΓYB��=c3����2�\gt*�uK7_��F?]�&/y��}���1��h��Do�+B@��l�P�j{?q�u ],)),���<����0��'�v�/�
p��e,��[L:ӂ�6�x.�$s��l�(>�H�i���+��mZ��
Q_�U��A�a���Y�`�!����ӻ&��7�r[�څ����xR��f��=aS�
�S"k{�|=���ja�3�m��ڂ�^Z3۔=�j���.��-�"�(�~�S��)7 ��|s�P=�P�&d��׸_�1�Kr�iy�KFB�o/{���4�5M2�z6���!��&����n)���<��.��t\����^~0i��@�N��:1W�;���3z�n_6�42�Ĝ�o� ����XbR�|�5�����eL�����uǰ�9
3��m��i�&P�8�2;�/c�-���h�̹�2ki ��@(!B���k����h8�qolJiiVm~QJ�h6_<Ⱦ��aZ�E���gw���qWH�$�4D��'��G�j �$є���U�&���򕄁�����D��Ilx	<K8O9%k��2�{LaM��uk�q�'���)�F�K#�%�Vë#5���f4K�Z����q���ۢ�`�؊i��[�/�Z5�5:9>�o���Nn^�ӳ����<Õ1��	��"�С9���k���lT(��� .7r�v�M�C!Fwy6��ʻ*o/5�-�Ai�ś�Ë��jp���:&���B�$:�iA+8d?���vMo��[�
?���4g�^wro�,3P[��^agu�W

q�v�(qg�T�1y\Q��.�����y���L�6����Fi�R�o��CJ!S��G!@����aX�����.�<1D�(/�	,|�´L��Q��i?�K�{|����e��p��Tu���T���A��ˇ�O9Q���Q�8�^oFu� |���~��-U�NpN�Y��YK�6yyg��� 5h�}*�*�6���Y�׭?F��ŗ���15�o@1Y����gfJ���t��8˕z�����^�/��G�U��5F�i5��kK�>�(�4� \��h���Y2ۅ_2�cx3�$���F�^#M�{+�\7⮚��39�~���p�F �H��=�nX��Q�`�E�F���*ދ��s5.���a��~+K@�1}��������$�y��^{��a~�+d&t܀����YA�}k.�}9y�d�J�Ue1���ph́���Թ�r%�u�<�{ˮ&,����7dT�\ӽ����{e���/���\8�Z����C��~z$ʓh�o�i��i�T�e2�͚�Ĕ��NRy�?j4&�8H�oQ��l��&>C>���r�WP`>7���i�Q�enG����������܈*����2�L`�gE�넛��C��s��_ e�7��^M�}B'�0|��ե�&=x�׵q%g9m�y���%>��4$ˋ�	��,�lT��p�����y;�<���,nω�$�&�C:�I!�Kۺ�u�� ����}v���n��A���9d�-'3q��4$���dZc�x6s�j�CHɍ�������~��!�D���ҎK�F}��m9�ˆ�ܜ���#��x`��xIy$w��/D"�M�h�l��#�|B5�^��}��.���>	Π�ivVz�+=p�)	`w��r��qVg�R������ݝ9���+��	@���_xw�w�+���)B�����p|bT�F�TSĐ��%�1֭g`?݌��a����X��W�J�{(���u��L��Ȣ�!�{l��*��������L�>YP�жF�g��w�?�W���I���<@A@��=γ�	�����[<�P@M�PV>���:3�L����>
	�s�gig���\�l���������|���f_����H�L���N��+�˲�#W��1�4v�t��4M�sZ�N|�>��z���&�a�S	�(�"mRn��ɰ�G9N�(���r���\X�e�l�I���qTfK�;���*�7��"D�90j��1p7��G8�ўg�-�~�t=�8�ǝ������+K>��BX�H�5�;���?~!oO~"���A=�K���R��ɜ�xn�m�aG��
�㺻:��$��
�+�i1m���=�C!�K����������i&d�\V�)yN @'���ҀeT
��oY#巼��`������Ϊ�<���n!6>i�3��.6L���o ��t��"hb͌h_

>>J�:L��c�O(/t�z}�
4:�`��
�Sկ<^�^L�?�X7�KN���CQK��ꗆe���1X6m�����(@"��oj���~;��j~����U�6fkLL��w�i�c	�+��S��E�Y���\V~Iqf��P =b���8w�1WC�:l���9:�eӻz��i�§~�n�ƭ�rU�:�.јB��'	F�ی_g��'�b�he����L���T4��4���Yo����gc��c ���^��r���]kϙ���@a_Kg *�&m���`��·aƽD�X�~0�?�]Bj��F�%�[�,��膄�@�BF�ȸ\ԧ��#�G�#��d	2�r8�Ŏʻ�d��Ѹ��{M�w�*�lC��Y��@��%Z��4�b�y."B���QGW�\�A��g�4�q0o#'ע���psi{����;�N��z��be�xˍ��I���i�W{>h�	���ܝ|	m�����ylr��i�_�y�t�,Zd�.�9�k��u��ނ*d��$����%�2�@�ɒ?E�Te��>��a*�T�U�i��2��djO$�����p�J^P���֮"�3(�_��ZBE����;���,���q`�M���u��g�H�Gd<|!":���� i��ٓ@�X�Q"TX�2���:������A
��\�-�ҋɡ�
�G��ND�� ����qA"�'gr�2=K�9��d`������/Z4�Ewd��m�X՞�b���>�]����9q���V�ݱ&� 6��4�u��,���LR�D��a}�����n�8�d���4n2�A�6�Z���d��Q�1��ʜ���4N�\�z�p;�iE�}�Y��
�ZW��j[���)��6Z���[�L�k$z�n��*#l���O�꺭����)�FV��}؟���{����p'��mK��#��V�
[��Ƭf�0ƔCU�~EȐ"ַ�����;ҡ���/n�����yA��P�?M��BjZCT��m��u��a��)`
H��w�-�z&��8�5Z���#,�)8��e�=��#&X��'T[hh$����G�w:a�,�hpަM#�?�9$P�x�:f�8�����+ b+L�q|=XB�UF��#8�-�q�z�����N�h�X$��'��p�-��~�r2"=�T=�AB�+���e4P�����ò]KMӶ[��>�1	D�`^  �B��
�e�Uo�Ԛ�|M���7���ٴ�m�\�~�$xk�����wpY\�:�C(\����<�SUu{�����d;rQ|�E�xl7�TDBL���1x]|�U�5<n�����7��y(V���+�kmp�Vkٛtm����Z�����x+l�M��'b� �@C�z,� ��-���Yt�R��7�뒜S.|v���U�V�lV���k�z�U����P�AKԝ,�Xn'YC+����D�9�U%k�	,����<��NH��hN̈�7O�ByK'�(P����j���pz�>c�M!���N���j�0�=����}N�:�OD�m�J����k�н�A\0�lYj�	�3��~���6K�$yetը��O�R7�i�z�W��c)_��=��I���+�#ήZ=��]0�Ş�[���P��i�>{xDZ\1��݂TQY����-< l� ����1y�6!���T���MJX�# �������h '�=������(;�H���6�@R�䑽}s��ғC�B�p��K�`�E�i�u��1v�gq��N�>V�Xs��Ǔ�C�������*���S�%``�E���L4��I�]1������-�7@k��8���C�'�L�p��AT���
���jfWi�Ov\�"~87�����:kݔɠ<X��~��ݟj�3Ke�J)-5$Ӡ&ś��=�(0;%����3���P	���"Jz��Ӕb�8���i{��6���v3+�BW8�F�П�,hU�����0x7�4��� v�'7F��}N}�@��W�? �j���6��-��f0�2Q�~� �-��\���b�|�P�^�����^�v�Q3,Ԧ]���P8;Q.��k��cXh�p�M9�(d!^OZ�\h�أ��\p��«'���x�D���آ}��_}�5�[�2]L>�FɶKOb�vo�
=��뙈�@��&>V�-�?̛~�VŷbU�ҿ\�C�`����"�ېjX�doۈ=:a��/X����G�<���p�p���������]bǾkM�o��!�}���� ӗj�PZ\�P��p����Io�	�|��#<8�9XI�S<\���� �D���$�Т���?`;��lT���2s8G�El�ͥ�9����Y��5A|�S�w_7{���ť���*zk��#�8FRKr\�l��$��. B�g�bH��_Ѭkj�M���7�]�)�Zd����a�C�-��h�C_�,�i��B��KCN�Z,����/�N��;Px!Z�����c�Q0�nI"~7��Z�����A�3��%L��	���V��c1y��{��ŵS�K0G5XQ4������l�ʁ@]�7�Y��
�3�ڔMj��#đ8�Jh���U�@�V�K�r��Q�H��`-�$'�y�	�1���lQm��g���Xh\~ET�X(�Eu���@��\D��`�VD޽J�s`n�E��-�~K�#eƋMe� EL�f��%`M�wv;��i^_�V����FVհ��־��%vG!o�K��vL��%c���a������Wy99��]N�%m��zڞl�*]R!x2��8��7f>�}��8�k�Ae����rRr8�
��W2L2�?�~�;�P���eT\w�]��I��lC �`}XN1R�|`��L*#GԨ�;�����(q�X�t���J��ș�t�D�6��n�ݑ�/�Z�AG�u-����x�Q3\�u���`�.Q�6�g< [S���c�rU�QfcO��s�~E,:����e:%ݶ��_Z��y;����������B�g�W��+���,@N-q�C��V��{���`�NS�TL�O�ݜ���0��C?��Mj���L��~yg�B/㓖a>��)���Y�h�F���x�.̛X6�Y�G���9,��L$����C���j$�+Q��Z��������@���l?�A	���{����7O F�/�~`aj_�-��I��Z�W����t�k�ʩ|�Nz�N�#,�����v�0��c��ccB�1J��@�<���<b����czMV6B��syz�?��٘�9�����<D��5.�I7���,�*t�l}��x	徸���Y���\�$r\]�⑰y76|;#��q��o8��V7V�6�>?(�Fp��C�v��d�G	FΉeT�W�+��u�M�����@<p@ �g�[���n�Q��uW��z���em>�'��s����N1/;a�؀�ڇ(3J�Y3Ca�tز�n�z�Yʏ8��[>j��s_�iO�V�=�`r$������5���jW�i��1�~���}�B`��MCfv����K���4JGq�y��6���Wz�Vd�ָ�Y4)/�پWJ��}L{�l�X]�e"��D,����zۃ|����-(ȃ�^?�Jtf����xg�w��L8	�9B�R��Xk��rB�rLb����aX�-��F��
b������Ț���L�tF�Tg@�J#��Y\J�-�<���U�ޣ�#{Y���
���v�
���xt��{J��1�=q��,�ؙ�M�a�@�|E2���M0i�4�^���4���Se�0���1��g�g��7~������F*��vP�4EZ?�Z�k�7o��t`C�6��_���(6� �8�4����>�`T(FNf�}��
�ް�ɝI�u0H�U��2%����g��ᒅã�8H��0�k$��Z�WP��W5h�.[R�9Uja@kBڈzʙX؅�&k-�Q�qŤL=,~�$-ep`t�]��g�vq��9w�є�l	UJ���9V�t��