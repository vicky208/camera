��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:���[�S�7�t1���TTI�[�g&�̍>�0�݁?n/��4v��O�댣·mjc��I���N@�Gj�G�����M��k��*�pcڑ7K�\7���y�nH��ab.�%��LѤx��u媠P�Xi�f��տ�S~
�A�O]�y����P1y������o��ғ��&�Ng��b�\�WN�nW�]�ha֝�ѡ�Wz�u�E�=bg�)3�ag2����֫��}z�hGgFѦ��!���k^��a�7�c�H�Na��+1�.�ct0���C/����y0��	Ӽק~�� [��E����]�����L��}!F��^���5��'���ZV�q0��n�����.:=�zFdv���A�T�>�w�''ꦢ�$�R� ���'j��@�²�*��<�Ԍ�l#ĥ(�1����	�7����Jq�]ul��h�X�|(GF����&�&�>)��"�x�N�U�����o�l<�Cho�B���8'�J�4�%jw4}xʠd�?�Xe�@�Еͨ�l ���@C�?����j0aBa_�z�����tϧ�����x꽰�Rّ/<�,�O�Qߏd!�%^V��y�}Ǉ�P��:��{��$d	C@%C����/��M*�3s��	��Ƈw�j2r���o��-_#!���
qF��t�V�;���hˈ���D���(q��wKI�a~s�5js��C��y�� $�v�=��_��h<[VV��&���f���;>o��P�hZi�o	�������0���]a�!_.��zHQ
x����D�w!z�K��Zi�@l�
Op����+j~!�(ٓ�6���l%�q�ɺ;Z��q)��T�Nf�2�����.�,��4�Gq�~�B���8(��Ｚ�	y.q���q�b|9���sM�j�Aj%�������%\�eY��vS�ot�Q(�!GhV�����Ԙ�A�U��~*�����P��>��:�����.3���K8v����i�u+1�B� �J_��hn�/5��*ݮ�!]���o���8�����K�<r�=@����+�S-6ܟq/���v=��T�w>.B[���3fHN@҇�46R��G#*%Ŕ,��)	-�Һ!����Rܕ�oBi��|�9U�́����������А�=��\~�	�?��8���=�)�[��ȶw'S�7]<њ`�f�Ơ֒����J�<)�r�+�
�]�r�dy�7�ʅ��x��}ȱ'|�1���-N$���2�X��l8��zr �{ʊu�])�Ư4�&��Rq͏4��іݭm��}���5v�g�::��.ǑA�����Azڶj��앣�	��س��)�j��M�?d��ݴɦXi�D��{3(��9��9�:-��o��[y8� m� ;]�F�1�W��5M]�OF�"�楁��3A}<;g5qq�r��� )i��gf��&��f�U-ϾD�;}�~P�.v/.קp�٩�E�܆��x :EY��.F�Ģ�����A��#�v�O;�&\���#�:��`��|�մe�l��
��x	k������qC�K��{��@ˏ�u����
9�P��%�Ŵ�0vݐaA�m�$��r`����G����q�nml�Y,Pv�u"s�)f{c�nܤ#Y�������k$^���d��� i�R8�����s�~_�mnx)��~l��/�
�D�a�"��[�RhD�z�����P��\�����q~	|їL�D�(���"�.�aT*����cL���Eb^|�ä9��
�q�,�}��e�7>���ޯ�
���[ ��ڗ���L2
_|���ȈP��*�mŶ�߱�&K�!z2?|�|�B�m2q!G�77�ެCR�D��gX݅�{�R�bI5 ���d���\�^��J@SC�DZ�vg^Ї׺j��#�F��~1h��Nx}��l�e�6�K�l��-�Yj�B� ��Kˊ%C��p���qk�l� t��V������]՗�%u/�<6	g��)4o�Z�m>89��z�'�y�C̿1��
�L�<�f���x��LսN�B����ŷ�Ɣr���Ę��C��WlW�*N�O^yȯύQ�V������^;�O�!Vg�~��u��|���wK�ZҦ���Ep&+�(��Pn����1�/k�H7	�y#����-���TYzN� p���?+��{�=��/I�>1΀FGgf\oI���*W��Z�����2���g�%���Y&ʁ���YPl�O�2��c�U�1��hR��K�
���k�(��֓��	�m�R�S
&�,��X��KV���A�jJM6��4��j�8���;Ne1Rq�N_���R{���:�h\RYIC����)SE�(]k�獌o�[��e)����p��c:��&6l۷��ZЁ)z�<��'uQ��m�5������Hj�O��E���b�Kh/T1=�;�&(�7
�XyzNv������z)n,R/�-��"�br�xX�zr��<\4�E�V�o8}:]csW�$`�����QpEc�#osXt�P���4�W;Sr�]�zn��G�;=a�Vdm&�U�#�I�P�4w<Xv�	6x�_ԧP�q<.PBJl;cW��0�C �Z��K6<69�"�;Y���.�6��,z��c!Ux�
h.��kL�5�~�M�hoŶ���Y*���#|R4Mf�jY�Xݹ^I�Ƨ#&���]t�O�8K߷֖�})��� ��J#�ٛC�5�!�T��.s��ASB�)V�3D\������Jk�?I���j*>E$!K���js����ߨ[8*�����i:Y�An�����-.n��z��L�f��q�.������H�i]��A�i���1QE'�T�AO=)���R_��3��-c��ͩˇG��;ykp��Γ;ǣ>]�l�Y�����t�v�g
���5��9E3�y������K��UYmѨ�1)�E0������̖��1�T1�,�l�S���������F��@AD�1k��J�'X8g��t��:n˟5kC���~����*�Qs��L�.�1��b���4�|��C�mTRݾ{4��� $�d�.��\Z\TK�,;ʟ]�N5��awp���($����{�9����9&�.��Z<(��;�Gz�E����֎`N��=�P+��H��v�v`�OɎՑ�R�����"���#I��~���<�M�v�q�O6�x{7�C�b�b�6w%���������W_dIa�O����L����2�"IH�=������c���TpƯ1�nYi���	�vfu��m�����/7��ls��>1���+8-(X|RQ�$��I�=�۪�������m�G����*)�u�q�(�ZJOY�-�e��!m u���ږv��d>ʼ�X���r0-=��J6p�0�{�ܔĂ �ÞB�Z��� ���6����ܔC���+ �d-�Z�z"�	Qڔ�=��T�)�ÀD*=����Od��`�t��`��)[K��2J��p����ר�6P�����gc�!���BG/��S�KgS�ԣ~��teٜ�cX���md��,�(�9e5���tx:����R��zk/0.�G�9$��c���{���.���S��_�fc�`��*`�
URX�j{���S�V�:4�>�4"
~3H������m�EȠ3�~�51)�~$-58���ɭ'@��<�N���?�4�b�a����U�SKY�u1,�
ma
�ǹ�py�y�K���HщZW���ML[�J���r�� w���sL�zE���8��Jp)�Q��!`�k�%��[���'t��֕��pe����Y������	@��>;峩 �=r'�AH�î��'���a=+�m���������]�|���Pm
�&.�E�r�bJ�/����>x�A���P�_���ã5V�wt��.����d�y)�ov�:���_��mh�v*�T�M��a�\_����^�?A���g��kW 7R���KeO��Ȼx��`��}�/���#	��r��9��\���j��c�1
h����+�B)�Z�<��%:E��#6Y�����f���!�d|ƴJ��rT+Ma�ʶp��a���4di�[��	HD���L��w���v>��F(݃z��qq���n����"���W���b�� ���fWӼD�K&Ք��J��E[V�@�]x�:Ц/fG�c�"��*��7T��i
tN;2���^�2�}i$��ģ��!�6��A� t���ߔ)9��xd��Vfm�Q�q�f/��+�o��N��
qd6f�`�EG�������%q��ۄ%�5�/Nvbj=!a�G��K��(�G�"h���z��ޢ�Fh�퐮���Q�nmeU\c�s�²e��ǈQ�Mi���+�ܼ1^���U��͐c'�H9<ۿG��>,��UD�BK�y�$2h"BeΌQ��8R��Bf�o�t!�ರ М��f$-N��C~}aRc�Y`�Z���~L�\�ǵ�#�-�� �����w*,�%Ʉ�t�^�ˍ]5�ie�C}�զT����%%��V9�j��|
*��~��X(:略���V��>�P锳P���q�m���6�7gF՗��gPK���w$5�qW�9����>(/�a4^��-B�6��F��&����Z�W��L�S����u �2IỿO�,�I��+@�Hm�D�|�!4!�2�RI�R_�D��sg8}ո����ږw���2���N����p��S�Kܝ&������� o�-Orۙ�&����NC�Ч �����;4��V�.9c����i윥�������*6`	����)�GN��:z�:_�z�:��ކ��xUA�Ȃ� '����(���ҫ	|�U>q�G��V:�|����d��N\E҈&�@k�C������T�4��d��N\���9�3�!d�C�"�?�^�ph�TÚ��i`���𲵅�(F �"�*�3�;lQ�L86z"��x����(v��k|hʙr���A�U�Y[j��r�ƈǽ2I��s۲��"`�`1�
���ӄ(V�X�0���v�T�piij]8qFVDY�6�MW�\����j��κ��)��ڇ+���q&�Lr~���چ��&$�(Ө�,yvn����n���\�c\ǋ��6?xԷ.%q�Q"X$rt�;�:��f��in#&�!�[J����7H�xA�jʙ�3���[|�K��)��'!:ou���cakn�(�_��`��uWЗ��v�E��Gt�0���Ӯ�\�nB���з�v&��S�6������H�g���T�[O��@��䖬�?�Ep�bͰ7�Td�,��Q�����,�o) [w�F̣Io��j��gG^M-���m�!8t�;Y�3�c.K_6Mw�˱���-9�pi`o�^�0�����U��&"U��hDZ*lD	M^}%�^(����t��k)P�Z�� ���f4�:�a�;h�-.�>Vu�䙤J�DSi��T���O�|ܖS��t5&k�x͵��NsĲ���9c*&�l�}��d�A��ׇ�^^ƺ�er�NF,~16�_������2 <ƕ�����uO�!�Ő���<$���?:�v?��څ�.#{�����\oSNN��Q���FR7�!0׮�R��R����6�)x[�z���ʦ*��5~f8L�Á��Sg$ͺ��,���;�{l��:[�]4x1_"�tD�	A�=/�+.�b�f�Fk�3�9�d�f2�ЍKC���1䉹5�����KPQ5wϘs G��X��Jn��Z2Y�g�t4C��ўf��Ui/���N3�m��8�0�P��7n" R'�2��b`�0����}�R����.k -	)���r��\j&h?�1뀲���!	�Yh���s�V�\"褘h�J0���|蓳�w���$�4�;.�{)�/��mC{x�3�4�U�	$͖e1ʆdS����)؃��zj
:�^���L@�<k{35aw(�ti� �l�`�e��ԝ�+}ذ4�Y��S�S�_���~:���0--|,CϾxc�V�,��������ȇ#��v �=�z!;%v��X+��tJ��Fx��x�_���C#L���́>n���ȡg�MVHĐ�)e/58y���t�6+!b��Aܸ;�����m�®�<�?��,��_�o�����O���$��pg�Z5>�t�R����j�0��r����6D8��}W�[��(�!��D���A�� �(�bmC��ID4�p���t����P��W�	#��癣�[N*D1��R������y��B���4 ���kN*���̫��2fO�&UN���fn=�+����ub�`�|l��ʵ+��δ����_�R�䫛�J��N���%$J��ߖVZx�nVI�����)�早�u�I�А����QT6�t�г
��7���ǹ�}��E�4D�3�{��U��R�ʔ��+���C��̛K`�J�o��OQ��e �.�x���g$�`���U����s��U7m����Q7 
��gc��F�`��p����!��k)��U��ywƖ�v8ī�^wt�}�yhò��(p�
���1S����|d�5	~�.22�8��	��TS���2�>	���3�wf�W�OL����q1�Q����!b4�F�+o��,���rڌO+���E��.k��TR��J��杝k��'��K�:՜�}�ly�Gz�n}�>R|�P�V�6'H�Z����t�Yմ;��ml&?����x�+�L_�h]Ƅ��/)Y��%�>�:��w����������g�7d��>�`�S�%�/B�� �AL6&��^!E�첮m.zt�'��k�jԷ���2�������hE�� �s���G$1
2T�����>��D)F��*�=�[��ha'���|�_b���ӡ��q�|=~s���|��IPj�t�A�`� �n���/��m�/�.�>k���+��KE�ly�=������|ZEAM�����Ԅ�6:&�&fӋC����1�����M,�����X��[�H
�+�Md��@*"Įء��M�%���$ny��F�`�:G;�+Ɉ�}E�X���}5�ҋ��J��uH�Y���^%{�{-.��/� ��
�6~I��3+Pa3"��a)u��L�@���o3�P�B��!�J��!�-&�D����ۻ��y׹}_S��*�n�>�-,�3X��*"i��쿢YjN���p�ؖ��J���:�[������N�8]"���q�~i��:�u�����c����/�l�L+�)`���?J�����H��o�$�WV�t�d,������E�?�R���:c�vBݺ���3�txzR�l}<��Ӛ�>�b*�i��iZ�FZ�󜇃�E��]&׎��)�B��7N��	6O��h���{o�-)~r`�Kui|k������|�-�z	�i/J��vb���& [8n:�����.�����(o��[���!�Z���]{��_�
���(�Ãd'G!I׬l%ෞP.N�^T�uՎd㚛��2x>�0�%?!)��aE�|p����/�J;��ir{��@�7TN�׺���-�2w�Ey��5��T���'Ui�����9,���$N�kw�G6�*��ޑ���YH�2Ļ��tss�1m�@��!+)�!8Rb���6վp8�N���a��M�K�o$�K�}�3_��U3�S�p�w� 7�d�� i����#��e@�j��Z��C��%��x
yc:�G���}?8�n��	�O�P/j�vU�q����t1�CX��
�+�5�t��*����7#Dl������Wz~~����4�i��pF�P����K*级D�ɗ2���.F`��	�u]MTrQ�?�*$��JuǬ(M� \#5JĚ�t����Ic�,�>~5~��ƽ��̧���4b,b�LIwklpY��+�-f����TIz?�{�u�\�N)�Bg��]�c	\Z�3z�W^�:!��,+� ��9wu���K@�m�<@��w��<����L{&�'�l状�*��(�իW�~��2�~��亮�#�<	���#�Zrb�/0)�d8�
���:;��� ��^��V���IV
`޶D˕���`׶�ӡ��Oќ� ��FH-���Bl��7(UG�b$M�k��*��8�l��ё�]�Ι/�W2ժ�5�X��U��Y�#Zbc4��^�z^�!D�!��2w�Q(���rIEZ܋ᇥ��F�a�Ӵ�n#�g�Ŵ��xf!�b����=�*�g�?����0c�,rǌ����cT�>T�BOp{�9�hrΩ�@N'4�؅!O��*祽�$8\�j�a������Pj��J�h\��F6ՙ�;�3̯�vD�逮;7g�C��EO����[ �D�a���a��i�Y����uGs*�䥦y��+�<4e�C�"�"L�֢'�Q�lޢ�U�����>-;�J�]�OD�$�v!P&z�Pj�=���X�HI�^��70���[�+����:�RB����1D[_3����N�)hL�?$�:!����}ؼ�ɗ�#e�?G9��K�/�ǋ׻m���&��
�������Z�:�뼨�v��*�y8��wr!EK~��]0e�^�ꔍƒ\�S��A��7]��Y��C�6_���}NJ=S�	�^�Rs���,�o|4wF��m���c��_�5��
��Ag ��w~���L��O��$9��Q�	���eJ�!kA�E
##��_YJ��l���-C�����v��@��zb�G�x�T@3�zch����T��y+n��l?���ޢ?��7΂�\�z����LGP��c�U�K���W��:D���:j$��6A?�7�Xs�������;�a��
����\���`7g�
�in>���D�ӉC����|Na��J�sG�@�����ؼ�8�t��MdGnߒ3�v������r��s�(e?x���²�lg�KW�; i�t�،t0�x1y��Fa�v����K�uG<t&��&4K4Ē�j��,J'Mˑfuݸ��~.3���X���!�G����=]�عfٱ̠.���T�!nZ���Ж�ao��H��K�:UY@N�c(�5�bUsi�I �d~T�}瓬#D����{�";�3�jn5]�(��X�977p��ztH���l��8S[,�ɦ¸-=;
6 �B�8�D+��G#A���I9Ao�yP6Wo�^���3�cJ�v,�Ǆ�\8Rڻ�a ���b�X$Z�`?���}�~؇��*/�[kwa�F�j��t _��v���3��e���*�?$sME�����+�d��7<Z���_�q�Jz�T�1�u.��3�$�:қ~����KN�,�1t�ؑ���3ŭ3bW����6o�уkƫ��M|C�	_wq�j��5�~8�9�a��e�}�.Z��*��S9_�����*��;_䧁I?W���j'a��o2/�w,W��>1"�w��>���տ���=B����C���b[�Q�Ӗ)�<�V��U\���-�&!��ò�+PG���'*� �����f�s�T�R��-9���������5�t�i���(��9=Q렓����l��`疷�h���C����b��}�+��=!��)����sI<�H��lg�n3��u�����{ֱ#��ad�b�Yw:9mސ�VMjd	���ns�B��ˇ?��'���F���Z �[���g�$�¯\b�Z�lW�cG-ݢ_�& �=Aݒi�ݠ��Ӵ&����,��p�m[1��,Y6�J���R9Į�zs�q�®U �FeN�C�|ɲ��,v�j��'Q���kMKм��N,��q9�9�}�,�2�����W&ױ�pR��V���;ܖoqW'��K��`\	pI
rl�W��0�"�@�8�B� ���>������t������;�e�o�6+���&ylT<�x�����܏�(����{*����$d�;)50�־��.U����|P?/鷯�L���%�K݆�?.�4v�0���$"�Rؽ@�i�� W�b%�#?Ʌ�Z^���g����L�9vU��%��5�[�F�� �z��<K$f��6���fʑ��&�t��8��Ӯ�A��kf�֤(k�UJ�y[�{�uǷ蜹����ֈ�;`��x������3�qT�=�*�#2= 0Ԭ+�C���kc�O��5ϧ�����k�= @5׼0�D3*�~�D�e2�~��ڇ�`�;��8�&6"gS����bjY�ʫ��?2��=]�T���f�1D�#cB����̔i��*�_t�[�����6����u��L�5���Z4�Ӓ��#!�!��QY�����w�w �`e�>��qHl4����m�\�*�!���U�D1 ������~d2|�c\��ί��䁚��o.2��6Pr� �,��Jl�Eѻ�w����Ǐ��RS%�K������a�fX�ɿZ�\v��*�%Iv�c����s��NK�$�@C�:B���(�.�q�i!\b�{�����4a		)"K�<��ѷˊ���A85x�/�ͣpS�P��*g X��w�q�`VS}���s�K ��a��y��na��=W� A�H1��p�Ǆ)��;uFԧ�K�v{*�d��� �_*�1��B��r��"wJgp�+66%�!���J GJ�?�4.�k.��%�rZcx�Y��g���UV��)ù�<"mxv~����8�P��;[N0I�Tz��''�#b J�#�f0J��1�6����~��+�.w��;HL�mgc����>�����R��y��9u��fٰ��V;�2T���Ac���\��(�f������Ԗ̯t�ωW�4X�6�
�m��mPyO �M_�`�M�8�uO�Dʑ�!����tU��
�U��K����t��U��s�V�z���βfvE{�A(5�$���=x�T�6�잼���ǇLN����M�t���I��e�НFr0�}��{<�a�mB�yv ��\����q2�2��Jdc�~ɺ�{c����g�;�C���"
���]���F�A�e	m��W�b�Ra�F!��yc�3|=�8�l(��L?�S�},(+X�7�t�B[mh,	vFؤ��O��������T�kޯ��|��^=\���`{���;k�u5�*�Gش�~�qWj�Ѷ��)���lk�C������.�E�Rl���~��2+$)�1�A� ���g:����j�&us�?��Vi��9��h�ۯ@����T�'��K�Mqk��)d�o��S��p�����r`B�=��e�ӷ��q(P�O�5����m���8�GT��#��D��(x��d�g�e�(e�{����a�7�Cy����Ύ��Gwc���6j����'�w�� 2࣢�<ud��FP�B|�8ӣ�a�]�UOv	��sҠ���럢!�҉,>#޶����g��Qv� �>̓,��|Y��I+*:k\0��s�%����a�vA��!�<��Ӝ�[�n��%��ծ3�K�C�E�+X8
X��d�Pԣ��?%I-">�g���*����}%�$A��mCC'��q����,��u����J�Y�GT���
`�v.����Ԃ�R�軥[�[|<���P1i/��9>-�"I]'�[+�iڐ�3TcʗU.9�T��W�?�6TiҮ�ϸ���N�-<5�g�mbS�'#��Nm�6,���0�݊Wf�'�s'6�ǎ��H]>����F�9�9b�1�2f����;�B�Q�Z��t�IY���M��$`pY��}�j�$ȅ*��UU^�!ζ����C+�F(}���Ỹ���L����X����dl����:��7��D��-:֌��s.Y�݊���4��}��K:���mITW�)x��?���_>��f���IbS��}�Ee떋�,����_�e�u�f{�/�����a���(�6���u���.�+����7���
e��p��׹!G�J�S����|�ؐ'7g�qo�?��G�> ��m��*n���q�q��Ne���}���c:@��� �=��ɤD��h/�1���4�b�V���Ԃ[=�ys����!C��)6Y1ħ0Y�R.�C��6dyTs�5~����`}�._x��)�O�W┟ae=2,'ܸ�R�a���u�g(�P�]��3mh}�;��ͣ���
YE��=��v+��@�|�׊�L�������-�n�ߢ�X��qs�q�Cva6���l��@��'#���0D3?��|_� ��2��Mj�[�^�;��w�6n���֕3�:�hE�r�Y�kԒΪJ��K{��L�n�4��wi�����nq����߼�� �@�?��:�Ͱ���:����4��E��u��Z��(=2PUR��{�_&��edBc�|��gnG����izN3��$X*�Q�L�����ɽD^��M�ՅJ�W���l��G��2��t�e�(����p���=u/��@.a��=�{��Nڭ1uK��5��9��
�aGtd�7N���pA)�'"Q���*�v���a�o|aA��a��i�Ӕ�or7��|�4g
t�Y�����: pMY����Me��8,�
�Ϛ;�����l٭$������J���w��c�%��N����X��+A����S*�@a��������� ��i͈�!4y2��n/����noL���cæ�nڰz�.~eW}|�W�h̳&D���#���������U	א�K\���w��1 M�5Ї�X�������xG	L�Z������4};��A����\���'�k;����u�f6t*�Utp��}��;ݓL��b{)���nr��i7��z�P�0���:zh���.�:yL������
�/�_���YA.]�T>uv:sq�D��SEP�Gn7`�{�l��tā|Q ��9��n��hR=w���l���7|�)��1<�<m9�[�VN�Ij޻/y=��H
4���T�[��MO�T�K��LľYu�hSM]:a�xq�:�ˑ{����M���g;�#(x)��I:w����k[��8�F��d�.����^3ȝ���>-6:lH�cx	��"oi�=�C��d�+�y���t�%�E=�|�/��aM�)��6 �Qa��>��{�Z�c������	c��h�F��}�ɦ�<c ����rS���9-�WeL�8���e?]X�kA��%c�,eY�YW���U]j���X��ߖ$\��ְ70��J������2��MHl�����*��w���:r�	�q&:�Dc�aB�?*�X��U��.Ꮩ�S�U�����Ä�dwp]�W�_���He�(�$wAL�
-�L�H{7�^��h��� �=
`@�x���}�˳H�ֶ�(�V�a��Z=��݆��O4��jc՞Ť�؃i����IC[MS��^�}d�H���\s�҈��T��(T��j�!���j��4�nYJ���5��Wh�^��"���4b0Y9�����Q�#0 Z�c���\�%�L.���$���8�c_d,qB�M�����_ā���Z�P�-x��*�	���<�_����Y���-�����bD�k�\�sg�O���G�e^@�Xb�t�����8V(ׅL�[�3@���s��;�I���%��(�a�k�:䶈�Θ�/���eΨr`^g�S!�����7"'�Y��%殦�E��'�d�*���U��kf5�I.u; /���2qe�ǋb��{���*���>��K��ѢE�r����WUlޛ�@��/5OX����%���B�Oqi���z�>��d
���c����:�W�:�(�8ӽ�G�φ�S�9/4?~��'F}���s�`�@���� HOd��'�������cb���x�����.s���� <�����4p���"H�Ti�#���.��(��g�7��:�c"-�?{��P_�O����|��|̉3|�
���C�r�	��<�_��J���	��	��&�9�a�?�˂�%�%d�F�*LBm��������V0BV���+�A��y��&Ku�l�͊�s�<uTb�4Q˷��j�64����D9��m*��1�]G�W�H�t5w��s`}�ŧN|~}[*}���s����5t��|���'P���џU��	�D�^ͧ	A���a�����tH��A������J�'@p c�Ԍ{ZC0u�ֽM�:��?�8���M*EJ-�J�H��J���+�I��6�%���
dr��is��]=�������3�
����EST�-O��T�S���-G.^`n��V"�+P}C��L�"o���-����D�=�:�a�<��S9֨N#ZG*�34x}��[��
�*�p���X�2t�.�ԉ�?�pzIsI�r�
R���~��]GU��1����݀�^�Ͼ�&�e�%���U\���*��K%l�6���DW��V�R��ZT���+?��=��?!a���2�>�P%�	#�����/�f�kՊS���<:�/ǖ7E�ͭ*!dK�Y���S�A-	��';Uɢ�-]���V�,�b�!���N�)b�����@@��F�e�Hָ:�ь�=h�������r�#c�]|���Q_���8h�� #�s�D��J��T4+�7ê7������ă��
f��Ȝ�v�^Z�AY��x��A���3�Z_9�k��Yg��$�q_��r�?׾���;�Fp����5l��7�Le�/ ��j��@a��� �Fj
 c�yh��*��;�ʚ=�܈7u`>T�0�X�s���񯲳�N"�����(P��*?��NW�q1�>�A�9�p�3\���`|x�S�cbr~Ί�|O�l��\{*x����_��&�g� ��%�
�x�B)�=�z/B�i>K�b��i�`Y��n������O24>�wW뀏7r�{Ѹ|H����,���~��c�B�L�*Tm�d��ұéhG�ò	�k�x�P�R�xa��B�x�)�Y�:�R՝ �37F�����T��[`��OEj>��ۭ0�$@��Vn�b;�]-NQ�r�E%)V��Q^P�wS)sk���bIx4�q"�Wa(�G����F�b
��=� ��/Vމ�E���p/:��2
�6���23�LX\�#��]h�q�r,�U�?�M|p.�z�_�Y�����2���o�� |Z*�J�&Ă˚�#��3ߞ4ư��*�C��8M�tS���M$����|c\�q��B�ؖT�,������]��R�8��Rjp,�T�=g��h��m;��A�
n�2o�:*oԦ�5!���$����`����jn�l��?Р���Roٙ�F�0��1�8�>�_�R�ѢPaZ�kd��n�N|���T�N+K�7>��j�x� ��8Hm�����'��(W������9S�!�� M�1`�6)o7�#�+�����_2�p�4gcH��X�۶E�.��pJ5hz�ɒx��;ZQ>�����ܜ���{��CGU��Zq��h��?��>\�Ņcô������*;`�5�Zg�)w�J����K~�&w6�.A@ɨa�fH[�\5(N��M����POM�G���%��?�w��������+��?�����2�&�p�:,�d�̗�id$`�-�x�\�}5`6G�i�p$9w��tyV�G� p����ya��7G_�0��T�v��"6��;Vq���.�>�#y�`�農�J2I9?�vx=��6mG ���4=�b^	���׺��MM[�}2� gf�y:݀ 3�ĦF�Z��P�Mz��}Y�b�r��X'��u���^ej��#vK�Z��3U����6�+����l{W8�f�C�Cq����[f �s���[嶏�$��_�z�Oi���F��q����7�1Z�N���_�������BaZ��|$���g|���_�q�{Fu�v{6���o�X�9�v�Hy*3�8��<���W"�����oø�qqqĲ~�)�"��%�<����^�F����C�ŉ���")�K�b��\ ��J�b��#�"&��gј����8QO���| ��$�H͙�Ϡ�A�<����H*I��Ek�W��A/�`�@}L��H~����\��4l�Q�?�G��&�im�U��[�#����� �B
/�s"�d�8��v||Uc�lW�u]|�K��x����j�	}$����49�ϸ��$�y����~"Pq�{�	����3҈�xS��7��{QC_�����l�~���3¯�!+�&�:S�0�aD#�p,�2�qj�x�Ƚ'Ԯ�
q5����v���7��a}^��Q=,v�=§M�t�]4	c�[ޛ)��|�B@�qN���tm�*�����AtGp	[�� ��J��7��c����=w�4������DB:]�p��+��l+]�b�W�J��6:��M)X9��B�t��x�X:�1N�X�1"��V�h=��^�K���g�=*�l�r�G�ȱ?�#����&]��ۼ���a��49���>�&>�L������C�e��̔u0UR��ߊ���pb �#����!{ �G��� �Wi��^����K�%:%�nX��>��4���;PSj�b�񡝠��۸�[��D5�P����&���a4����	�!��-�;�w]vcN�
ZN�ǋ��q�yI�����E���c��A�F����T}��`[���"�-�+��> 7}����ZF{�{�r��;u;��PK%��4?�Ve�F��`6t�#u�X�� ,�{��*�]|Gg�%桚E��xإ?է� e�qӱ�3^�O����N�zGEj<�3	�{��+e��������� Z^��x�heV���Z�߅u��T���fyi]\�Mc�f����Q��CK.���0�E���b��#��t�ٔ�\���,ޓ�B��y��\:��<�^\�C�R�̥��l�b�Kۣ�4a��K��ef���ƑΝ��b�?$!J�V%5�?ٞ����	�>������!+]� ��>���6�yi^�>11��� <Ge�>\����������0���]��F�br4`b_�={�'�E�P��2l�Y�N�2�|c"W:+����:��#���y���N�o��J�@��:�:�~�dKӹ�����
�F+Ws�ϑ�4���2;ѯ��h���aҪ�W�P+h��6��i{r)�J�%�Nu���e=֞�\x��������U�J��+�%_���M��+���s��X�}�?�j{2M�y�`�<�+���$ ��?k
�tSL�re����q�&5�����Cd�V��h����zӜ��3�����2/�wH�J@�i�e]Q_s6er�ѕ#JX�9�"Q�5p�5�C眛���AI!�Gƺ�99�2�!p�eP32d+�J<v&R��G'��zC�|���k�����D�}q��%�C@낐[�<Յ�-c-�A���uU��"�us�~L�0v>���H�j� ��.���F��{$(,�;D�>Ʀ�A��Գ�zG�4���S���n��C�$*u<��ܗ3Y���������܌���lG��	��
���D����N5\1�������7���}������Թ�{�K�7w��t�����׸o�H �*��-E;]ߞ-4Z�����e=9��*�EyV�[3�SP׫����7���~tZ���#�5i.o�@./A�S�IXMub��\y!����M�=f7�!���|�?̬ k/t��J	�楬�}�6�Z����gyM�:��!�WAgG+u�&��L�q83KG��dQ����#�)Ngz���(�L�Yy��֚��7Ø�U����&�Z	�;@Z�����W1��<�8sv>�AX����E,$-��ܧ�5��u��x����	��Bp���K�'�t�k#��K'ԋ@� ?��*��^��Vk����$X�%���2�(��ɸ�OC��e	�L�ojQ���1�.�<k��֍N���U�U�<B�d(�:k�ݚ����A��D_��.4�������=���ra�O,���a%bO���'znV��nTO�㌩S�*y���v,�٥WQ#�P�P�����X�4����BCM�j"�-Oh%�Yޟk]�l��V����/�>{Y�S�&i��D�b�bڶ�kʤ�m�,	�Ջ(�uFE*r�N�iv�7���(��Y[��ca0�n��\���DD�䰠��ɣ5�5���"�9%.ǣ���#�����]e.�����f��VY��iR��v���E��e[=%����pbֿ>^m��v��5���$��#�FW���w�p�*?�g���˫�~}�}�1Q�!��\:'��a��/� Dj����sqv�M<�/l�oZ ��*sG�T��m�af��Q���Ͳg�����M��s��e�I�OE%8F�n)n>n{� �PH��{�����g�n�&n�i��Y{�k<�{US�y��!s&�u}�+��A����p�դ��^���ihL��R�I��S�O�Z�y�w��<�p&��H�I��M�s\�Y?VC���U���!������<����e6�{1�/���a14J���̪������{XAG%���N0�d
�Ƕ;�������!���bͼ�q��aK�֩�7�?,B�<�2���$�Y�c�2	�S��L�zE5��9PM
7A���m�2���G���wE]� ƶt���Tͱ�g@�
���3��;�\�lUE�nH�"���Q�jbP�nآ����;���w�v=}	��k�M�x�Ҽ��I�����ߧ�P�3�%�r�|��f�I� ��^�����6���HC��7K��v8��K��r��7��MHN5�ޤ�8ԝ3
P���*�L�I\��
b`�!P�|��i#��Ru16����x�K�)`t�v�P]#�(	��r����/�(�����9�P�W�]p)��d�Q�@tr~b�+�T�ڡ.Dǖ�f���3 ��ˮ��JjX��e��a ���P�'W�_^����1j�����;MX������w[�� � �\Cܢ z6�����n�µ�"�(%#7�=6���oSZ	Y�8jE�Zyd�:D�H��D%W)Ib}�}w��J��O�"~�5����J���R���$|s��R�RXM6u���g⩑��;�j��sU)K���c���jМ)�H�4�lEt��`\w���z즍0M%Jv�H�����\b4$����qGh;�ڏS~��&�h�Q��序�D�ʺ�/#�u7�n7ו��D�P�S�<7z8=��T|�.ɱP,�M[>�!��������󲐒F��$j��+�]�ۘ풦8J�5V [�K�H��r*�����$�	p��L��@ش��|�+D��2�V�����|Wx"�K@Е����ʡ�F��ή�+Yx#
	x�����©T���~
��d�����]av-�����?�y�5N�x���|�¸��xqT�h,I�~s�fhL��y1����G'�F��C����m"Q�� ���������:%��B�`���B��ꓝ/H�#;�5��F��vֺ����:�Ea��Oٸ��G�< {_ˢ�h��"�o�=)�*1� ��D@a�T@j�dO�F�xm��<�^�c�^���9�[�-�@�˿#T�����G�>.� /�\�)�s���0��<)$�tS�J�Ag��U��P#��#�;��ޗ��ss��Ccdv��`�8}�%jm���2�{éS?��7�HylF���.5_~#GFOy
k��x���3�k)���o���FU�����fc�V�S�Tw�zE�e7�o��J���'?J�m�;�5���(����#N�قS_��X&��x�;�����pQ��K��~:,�N�K���m�Ӯ���٧��p�&�S��l��D5HDg�ֺ�uWC5bb���Uk�)y��y��/-�xZu��ca��
��|��<�S��d���?�អ78C�n����R&X��J8�� ����S����%a�=J��;���Y���2Ɯ6�s	����dL�=!�vp�4Cǝ� ,̅�A19�B3�〶�0|[��w�A���c�W�~���2� u�=)����1Z,(i�19&�!��3��'pC|8M�Vm��e��<*w�B�Ɉ� :��NFwr���޸K7������B�-��J��{qOڵ��~����7뚶~�w����cAc�C]2)�����@��c�� &75�L��]ѩ+�-)���52��	(F�R�y�Q��}��b{�Cf����x<��s��)Dz1#=���hhȗa���PJ��D���@��؎�?�{�k��eH������=2c�aDՄw����c��UQ���X�U'��-�KD��-C��Q_��<���7)j�|`��8Dh(C�O9�Ȟ �
l�";��$��
�У�eĕ�vȃ64k�6��f�?��8��n�=��s�f�����Br8J��"e�X��F������W/x+l>2��S��IX��m��P˔*hd
�h�����	��\�C��	��ZBwʟ$�	:$L{��\��҈g�Q��r���7\��t*M`h�Y�+o��5��F�v��j���S��N��i��@���q�2�\y�K�����d��l]��֙�5����Ez'��CKl̝�ن���7������k)af��rp3��4c�l�a���kD��a���TD��� �0��)�cI�4�R��L/�JI�iL�B�O���m��j�(ⴼD)�Y<���@a�t+W7?��x���]��w�c� ��M�����$Ij^��4�|8���3��G�9���R�/B�g��Q�*\H�Ʒ49~�����	��+��
o2PM&:����W�3�I�G�rNեMg��:C��Ov��^D"e�p���p��O�P.�nk֑��>�n���?��0�V�|����Ę��G�4`drUk�w�	�a���7��}�1pdD�|u�G�Cx��EGE�o�&�o��`�p�h0c�Ӻ�(��#C���R���	��x������C�وk����q¿��}(�1�ٰ�5ڗb�	+��P_�Z��[�Z��(�����t��ã��Dv*�j�X���
��1rT�xX�ܾ�S7�Q��р*֌]؉a�1<s8]\m�g}�|���"0Vh��TSq����ll��'.�/.]�h��:0����4)���Kx&�.�ò������B?0o��7y�9�U�ᑢ`rX%c$B�*�'>��������P�� 9�R���� �j6�0?ڶ�JѬ�큵6���P��Z/"jU��q�UZ��q�gi}rq���R&�
�eq깵4�bqy
�٧�����}���jd92{��� T�Y �ZペD#v2��ZDW�j��s�,�r�Xe�D�\u���S>Av��Ukcz�	"�.[͐U�A�_�O��_[�yC��#��:��k'Zv�B듼V� (H��p��;�b*0\��[ n	ю���_e�T���`P���'mI��@V5�L1M��7�Ȉ����֏s�M�8��+ª����E��BR���L`�F<�{��6Ϙ!������-��޼,b�d�t�ϻg_���yoW`��s��(պ*�j��T����m{*]d��u�W�����Ք��0��Ư}4yY�w��o,w+_)iSÒ:$�?�����gF��i��00m4�˥�F$w���FOʻJ��N�J=�Y��щ�3Ƶ�Ў3mH3�H;�Y�X'���Q��t�ڣ��J�r���L��	�^ƥ�
%�ED�l�%�I\�L9;{�<m0�4��3	͎P�^S+��4K�*J�خ0��jʹR"�LJ;F^�5?�|ba~q�� ��RR�X�;wq�^v�}*�>�OIfx�Ŀ�v<:�_1m]�4q����3o��F������u����)�2e*ꩫ��zp}ܬ*�Q���`8U�E���a�З��
��s�j\"��[�<�!J�͢����=9���~T�P�(��	W
�⍘�%U���<�ml���O�i�d�i~c�*`B�c����"��z_s�]��GZoDa��m.}>��u
^2���'	3��q��ŭf]C���J����$�����I�3�-T�R�p�e��|�|�V�lfpD7�y gF�,�_�!��M�)��d���2���&UvV.cx�Դ�-�`��@��G=kuF��qE��gcx"3H�X��$�z\�'�2C?�f�kyw�nQa�����
�X@]W���,l��	�vqN3�rH�מts�;o��AWX��d���:��+<{a@d����z�rG�>�W�g���D�yw��7M��0� 'd��nK����V�@em܇���Rvl�P�HA�p1���k�'cx �Z}����G+5��I��99מ�w'�P� ��!M�Wh�Zh2�[>K��I������3l��G��_��̝N..$\_�&��@������:�$����+�B>Z�0X�<�;�Ӵ3
��Fo���z�(0����Z��6Q_*��!غz|n�#>��1�v|�&�o�hٰzBV�)1����r�ub�<8b�먀��c�rv�ט'���E��k�k�49M c̓��J���%�M*�Q��k�9��$>�$��B�B���ѮjOrE�e��z3kS"�9�9"I�&n�"g(�+�F54);QP�8�gA��"K�1Qijs駛<�!�|����4R�@k�X\�(��GS���Fa�q����J�uw���WT�;k/���@s7�m3�t�� �Ms;,�?������r��@]���N6֯����k���O�K������9�`�O�u��-Eh�#jHO�RIq�,>�hZ8>��*=�*�$�gȷ�d��5����<���"D����6�R�������?�&�7�(]M�岹�nJ�Е,����H�T�;X���2Za�iOC�q�;|�>�ÒW���.�4�L������N�I{�J�r�D�x��9ٽ/��dOc��v�kP�413�Ӽ9�w������0�.��*�u�a�_[��}@t� ϙ$���qP����s��;��t��a٨~�j��v����	X�U�%�q?ݳ1.��
~�c��1�����0Ab0�9��"bf�����E��߉KqE1p���~�����9z��f�K^���*��9R��0�]w;:u�
gנ�r��L��w7i����7�xثD4�$oo��`��jh(Ћ��%� u�u|еu�e
����&ΪO@�GHu<̫�V	�x�pt�0�9�c�r����PL(�X[�vR��5W�:qPia��u�8r�"��ePfn)8��P(4O5k�A� Ó]�h&�('� ��'w5�3�A��u�8Ņi��L\��&n7�,�.�)��H9���|�k��K��U'�L�)?����w�b;��l8�"����d��i�/<G��d���S�ԃ.+�b��2D���:g@��Y�l�m>.e�p��*�rj��.��)��x_s��AK�`�P�E&�^֕�G��ZX��^_57X�!�ix�b��y�P�D�L8N��U��:`j��l�/��c��>w���	�����M��c�p�k��FP6z�1V�B�����Lk�E�N����Z>G�y�bQ<��m]�8@�WTzu$��,��C��*$t����]��~��QJ��P���	h��H:)+�5�����u���%��P
�q���y�V�/��>�|Oӝ��x��~d�R8h��Ta,B�\o(�
s�r.(-6mԄ����~:ӭ
�-�XƏ"^V��g�Q�t:�Ԙ��`w|^V'V�9볬��ᾫ��u����=l鶴o�H����0�K�-=�G�L ����g�={�����I���IE݀���x�^ZW[�D��D��+�6(	�5˚+���n�U�"���!����6�e �N`ӸM���Q�y��"$�_8U�]�qDg��b>�7|7hՒ�y��V����B�5�4�/�/��
/�E�TpS��4��F��E �W���9ߧ�rR�Mcє|Vݠ�v���s����z��C-B6-xbUBqUEpE� ��y�~�i>j��J���������p��YLR��r�X�0�>������n�R��D2�I�h�3�X�͈q��*#c#ѹ�4��Xʙ��ut/�Y��M;}��	]b�F���?�}KUԍ^߫H�;��m���u�{����Ն�L{,�~��V������D>0����ì�"���A���� �vk��N�C�SU�^�[���҆��+��5��z!L���0��՚�������I3��IG��}�����믻?���U��O̓wK;�^֞�6�u�u���,�W�E��tcN����1�ˤ/s�جZ�E�jx�cXڧ�H6br��+��{��WF�C���O���B�V�����&��Bǡ�m�Q���1��s�*(�)�9G�
�%���4k���Ͼ����7�j�:?���V#���&��}�ܺ8ǈ����-d���U`v�rjq3��bS1�F�����޺��y@P%0'ո���HTa�D���&�#U��D�:�����\U}������y��/�BK���j��$��^����ozz;W߹xa�#R���(W],{� �F����M�Y���Y�5G3��9R�2v)g��4)Ƽo�g�9o�-�'E���-�����0��,R��Ltُ��n�I���?{�]�ʥg �R��b���8�Z8+V�s���$����!��C��c�
=�m�3�7�-�#�ҍ�z�h���VSa�BB�/3�劏�����n���T*=̢jL��@�0:�HD��6Wl&��r��Bt�u���Y\�s���?�xj��CZK�vkS�3�4��g��F�9�덚[�o �n2�z�Ъ:)������
?��ў?�Q��2�[Ф�96�e�c��=p�J'� f��G:7�%\���W?6{g���N����LՏ{7���C��gKKs	��-@j��A����GIx�_�X���W���U*&D�_�:k)�}��^�񮎘n�pu%fG�-�_
`�� u"�8�	�K���X��p�y��'.B�LtM��}GjZ��չ�H2����~�_ӥ%�Y��É���^}c�
M�Q�˕.$�ɬ@�ذ�9n��!)^��d��+540�aw޳̚]���',WI�H���?�������
���TƆ9��_��_~�C�Z�/�������,>u���lT��½�V���
sM�0�gTQXΖ)*��) �M�*<����	���p�"���\��S��;�H���To�1ծ�?��~���y��D���G�+E_xG"@M/���E�vW���ᗨ�Y� ����/�lm`�Ӛ`�c�
Z�|e{�v�7�J��H6۾|�W�H�t D��$Zּa���Gwr���mƇ���i�3����Z.ee+�%�٦�{׻�n�����"�h6Ͷ��1$el�����=nN����I���Nޢ,��>��v���05�d��~�_�XKƠY#Q�iс� �T���kQ5�;_�*���Ik	�ɼc���_�
_�3�̮���ڮ��|D����%b�C�[
��\ga�N:�I�)b:2_w�"�����܎�����v��SCґ/Q�@���n�mE��m�X����ou�����"�@�b�Pq����M��8;Л�9'�����gF����u��jt�V���-CR�sD5
N�w�
+xU0K�*�l��x��l>�Kv0v���p��:��9T�j6�P�^Q{lf�_�|�>�ٸ�1�jiv�ʾ;����D�9]��o����x8T2�e ��Q���rn.~�-֦��cҏ����*]염���U���z��zԥ.����L�S8���8�<J8�κ^jy��~�)=G:��������ыp��٢��G��Qg8�7\Դ:J�g�ޠ��8���V@KTmA)�
ƱBb�:���Ǌg��J>�T�����#_D�=�z���r_4,Jƭ�A�������؝]��3��7�^���+x�d��Լ�+!��pϠ�K�F��.��8������ʥ���+�g���_�		�l�B����7Rj�X=7����hLBe��]ϭ6�=�p`>=���ZA�QDY؇�߲����`�`7�_�I����m��0{��;�QXyD�
��;�E[�o�On� H��S]]R)�,a',�p4��>�����=���I��0��/�؊�p���B�UH���u7�7̇�i�6�3��i�Xj�z2%����D�=.���"�Մ�l�;���٢/�i�E�",	i���J�D~����m<-�!j�H)ef.���7]hP��hև<Ra�1���Υ�Y;���	�3+�,�l�*��KN�IO7�qBB�JS|�!�Ǡ����oh����3��R�tT�V;��Y8�xaLfRQos��խ�6��nK^В���(c�d�/�R_�|,h7���V�މg~��H�W�IO.��h�J�˴�Y�O	1n�.�x"��T�t�x˿�c��l���3n,%��VT�hO�Zf��!G ��HkJ<�v#&��v�ޟʨS$��p�����k�ԉ���`}�0�ҡH�7��z	�Ȗ0I�o�N~��IVp��$?����a�u�e ���}��ظ��7���I���X!1ikH��$֯�o��KW�K���&�Op�`��p��r�D[�(*�ڞa����n��j��yZ�_��'b�:���(����M#/�$˜�
N�_H�3��#��Qb>�?(u�0�p�sn�"��d�ކ)�-��<�����:�r|]�\�GÉJ���9���eL���	��/Tw�?��$��pL�1�`x$��Iܔ�a瘑]kදW�q��k�r���"[����^ã0���;�?�6`����}�Q���9*��d����S��E�Su������Iu{���9�}�N+A�C��x"������3���v��b�Ec�@t}�z�{m#�pS �i6��ܿ��D:c����+�AY��:��\��;�i)PS��L�V��BA����c��,ۯ����E�g�>��,�K�~���mw���tvv�k�^5�bƫ�{�֧'g�}|�鯞�?�D����S�(�kgq�^.�xॠ<��[-�x��$�bʼ�%�����N��zf�i�x݄�|C��w��S9j���z���7a�'����~�@I`ȳs~��6X�Nt�dL�UZ���R�����c��5P#�,�K�'���m�5��1D���(�n����r��'x�gx;�{L����u!#t���$�1�t��!������t��@�mWz��u��;���N`��xb�Z���@Ɠw�J�WI7�����1�5��w�u*���S��;����]h���?���c���nw�[��kx��,�ۨ�"�!9����;������hEN�S �π{9��
2�s=�8�8��K���������v�ޢd�4��7H�I�@��*�$��C�!��L�ax��~��Տ����.����.%I��\�����"�u���z�Barr�)�PT^�!����H���G��,FbR2��f
�����'@|�cu�6Ta�c7�-�uq���7�'e<ԅB'Ȥu*�͚}���Fg-�v��'P2}�cDA��ґu��X��~��"�1h̴�O$г0�O����������~U͇m�:P�&n͛^	IH�tv�-�՚ �n��\/����2�+^�Gk�YKʬ�0�X��C��![Rx�Q����A\xĩSf?�C�ᕋ/#Y�=6C�}.�T�o����������e�1��tj��e3��l��P��pb�J��X�Nb6X(-l݀��Ȍ���(�<�W1�T�!�h���$�9�x��tU��b|?�,]<�-��^t8qvF���]x��ck�FV�5^�)��^�t
	��O��HX�ʭ�(&-�ޝ�6�ծ�$}0c���jѭﵽ����a�>��Qt?��}^m �v� � %!��f���bM&%gA?%�n��;������4�I�7���!v�̯֭7�F���,�"����J�BQ��&�.Vm�l\�q�?���|��q;Z&T�Z��:1������j��� QA�vg�/���4%�쪃źL��v��'PB�25�o����5W,"�lR��3s�_Ĵ�J�Y���-�U��Mp�B�8'�ˋ�8���m%��$������
���J�ݮS�-7Q�z-_lp��B�!��Ogx�~�@�C���}dv)����$1���0�Ԭ�S�֔��A�W9N��O����6�N̋�&�^x�B.P.fb >��L���O�TE��&(�F��	�t4�,և�t��Z�h�������d���
Ĵ�ڣJՋ�	&�hx�-�ߏw���8`���u�(�_u��xct��?�pEh��镡�������bCx�36�!��'�7��@`�F�$/Ҹ�i,�b��m��p��y#p����ݩy_�5�n ���*=��6�J:\��j>����{� �nŜ3���Lʰ% �9�r�t��v���j��x�"��}����\�o^X���̨\�\0dٲӢ7x�}�e-�v4n'�C��Ԏl/��8V��/,+��K�6�Ԗ��"��
HwKSS�9ܵ��w�Nx�*���v<����p3��COPNv��!d��� @�k��T�7^���E�g7��Ff5� �?ĕ���N o�&��� K	������@`>0}"�$����*�A��6#{���E~�q�%���4��xL�n��C�8�M�	�UP�*�Y���#���v;1J�Gq]�:�;r�Lp�o ��]�ߥ�d:�������3����<�P%#�3.��A��U���"��&����	�=�~D��ij��\[�?E�(��G6��8K�F�w-�I���t�F�v���)dzAUsTb��b.ŲaXV�х}n�B}���Ю�f��O�}�Q����b�?_KpL������� ��KO���$@�"J��)V]$��+�67�ʔOh����v��B>�?��%�U�/S�|"�9���n���Ըwv�P|"�9qCU./�Gw|��N"b��b��u�}���<�ȵɚ3ע؛�"�]�@��{>|<�³��ޚ:�xt�����~���W ��S�]]�9��WY:,��P�˚C0��&�=D��f)�L�Z0%�����<'o���38���� & Hڄ7$�lC����܍6}B��3�o�2�ë�3�'tJ���`����a�]�y�NƠ�h@�*��T�� ����wf��fa"��ɎS$������i/���R��k�Y{'e���N��!6`�mpW?1�T��E�B��#�D�'7��,�-q`Z�e�7�����A�.��g��d.zc~�k	�}���h9�	ߚ�8�D�{�#��$\���b�	�iP����F���|�5d��l�'nj��lf�h�]�w���F�Hꛗ�k�7I����Z�B��,�t$*+Lm��G�S������3A)Uq��Z�O� �3��`ZJ�^����obl���g�Դ���,NXz��Nϒ�w'�>�P�OZ2�T��/�@�]�Դ�����Zɯ��wݗ^��)�;�l��ނ���h�^jbXmL���&�Vh�H���]���げ��ߐ0�.3��0�8�m��q��ش�i�8�
���ͭ����́^%ȿ�/D�m�LE�W�j��\�հ�������j[xJW�m^��H����Y�Ѳ<N-����V0"��U�-�o#i����o.�U1��%��%o^U�-�.��q8�\����H����ߓ5?9�M�@֪��Ƣ2M�1'���S�
�B�|
�w�L��p"miXg�Ƀ�!�k��X����S��u��t��k~o
�W��J�1�B\{�K>��J!����#5hQ����22�{ �me��["g��7O�j@\������ %P��⚰�2���E\�O���Mh��C*7jU~�����S�0T���ͣ��������$���RQ��V�J�gQe�(_O�$�Y�z�lOІ����{���I��C�Vƫ,�6�����FH�n����D�&.���@=��%p�1B�;����}Lm*���ݨf]B�Հg#�W��ѭ}��}��~����M������qr-q�O�q�<o,}Ԋ3?�@4J��a	`����|�l��H�V6�Q�<$�+Ώ�5eK�}��S+x��݇_w��_���O��1=	�~��[�eS�&E���V�Ź�}J��A��+�'ab@<�8����3~k����V�:i ��~A��Tb�LF-�#	�F�d�Y�9�O3��i�nw�?��ܱ�r�0�mG|�\j;�m"^���i��g4���x�=}���J ��kz�$��t�OG�,�@�􉧎���t%=��ִq����ۍ�c���*s�K�p����<�0x#�ҧ"�1` T��h��P����:�V(��oCF��%��)�rM�駄��]�VLA�jcQZa��N��6*����zrQw�\�$'��q|P����b�ht�M��i�n�]w���b2�7}S�-���p�D�"x�~E�};�%�[�����3[=}�D��v��C����X�>F{��[����7A�Z��7�@����x��6��ր;;��Q?�̔Q�ӁׇZ����������~���Uu4�Ο(�
j��`�w�k���)i�T��x�}ڰ�ұ��6�ĂC\D�p�׫dP%��G��O�xԚ��ˀ���:l��ǣ�D��h�@N��k���s��Ϙ�@D��������$�/Qm���A�p����W=u�]9÷l �l_\�.U����^gkH�+�$��sr�HWނ���:`w��$��hx$x��UG�X2K�;#η.��DjfVk�N+Hx4���߆v�SITЗ���9+\�~{�f?��D�j���gl6��K�űmS�!&&�3I���Ԛ�1^j����ݧ��ƣ\`7�]��t������ՑυQ|Z	Bq9�C����Z��{�@0H.�C�Q8���?�)_N�Q	���Mq\��}�u5#�=��4�J���b�gc��0����:�1��o�݈�ds�fDȡ[�B��(WTZ"����qqt�ڽ����'P@���f	@tl�c	����k��}�v�b��H_T��7o�7��5�-97� М��gL*���q �>!�툠��(�yI����N��@Oǔ���w�7?D�X�Ζ�����+ɒ��I�f�P�7�xv�E&1�	iu��dc���A��$�UȚ$��)�J��9��ů?-(�]JR�!���ҕ'����鰖�1S����Gi�M�T�U6G��+]\��D���HI��
��U��?�ԤY'�d�r�ב�d��b�
�nhq�<�alFc�������%�Ʋ�(��9�1��Kf�C�A�Kv��/!�F���V�)gG�a�+>�%*�du+����[��tmA�)27�����Q���H�,��_�D�
����?�Q��s��#���.aģV���}Y`��z�����h����Uw�r=/-ؒ��q��q�k�'t��K�j_�1綪�^8����e�����it�}���5�Z}��Vqn�?�]�Q����S/�����{[$�g�'�Qf�6�I�k�
e>c7�����\[!2{�I$� &����*_�Ƥ�4���>4q0��~�4*��N7@�&��>/s���$�i �%;g���t�y�م�7�-��}l*h�d��I��)ͫM��JzJ���h�gDX�"��#�&��'� ��^��>�l�
�oo�{���L�_����G���M�?*�W$_�Mܫ�T���2UF��l�(<I��i���K4�_�m����&�yŚ+'B�m�_�������D'�
2Pͦ��v� "�
��!2�.���H�@S�6m�%
8X�Ȟ���t]��t�MEZP,����K��rY�k��W�ʘ��A(� �̧"�=-(O[]	�/?jSM�oM�����8������@����9~�
!�Z$)��֙n?Ú�Խ���U,u�ܝ�Ě�f���QdSG����\*��Ӓ�Naģ,<+"���C�K���B7;��a��51���j�RK�q��ֲ�ꟴ?�L	s�=�h@B�K�e��ᆘ.�h�{1�m�4���t�i��Ʌ���.����^��[�k�r(��[8j���n��Z3����ߋ�:}0G9�28`Н�Jɘ�Q9A�ĭ+�����-8r��gk�s�u�����r'�W$��9c��:�U��걣邰 ��g����ܹ9� �Yy[��x��V�&�]/_U��r�䙬FIk�Ӻ}�>�׹���dJSkE�
쎭xϯ�t�9M1?�i��2KxEP ��a��H�wv��;��e�f2O�+������˝�4G�.�\|�s���=
��ȈX}~���L�tߊr;`x�,$s��H��-�W��w���K���x,�
-97�C�8�&������.� @z�e����w�����9�h�D�̟�r��>�+g�s#?�'���>���|����zh'2"�����c����]��R�X��Y����f�P��������z�N(u ,=�D���%��K�D�֩�ߊ�A��`>�gڍ꜉e��"��+//�0���y33��#wo�e��ޑ��v�m��<2�|���V�z������ ׁ��QK/N��}2�@vEo�B��ed{T�d�7/O
	�=�!)���g�T�	��5e�z��4�A4߄���k����E:;��_^\?�ț�"��]e%���<u�9U5(�"�i�u�\����c�DgGP]�!�
��4@T���χ��id<�ڐ��vI�[��>�d�W6�o��E$%���j�3����4oK�6�N����/�=���}�g|<�.�cʆ��88\'Z�`>N�#�7�׈��oД|}͑��G�[�b����mhs����?�]D�ܭ9$���f�B�t�C�S�+�yF�h0�f#D��J�Xb�gX�*{�����:&��:�FP8஀��L�7l���fB�Q�����T��v����nF��X���v=�xП�ʭ/�zQnP���^Y����YS&��1�A�s���ܷ)�a��<P�/S^z�s��?� �����XĊ��9F���I
`��c����;�{ٰy�y��d��&*��V���ZCGW���B\���ۯ ����K�-���DF.�ì3&!^B���?��@C"~�.����n}����[Y�c�3�uHr��DQ{�D�E\���������&ߓ�@�i'�3�҉��e�YI��^?�q�I�^3�z�>2�y�n�������������o�&�;9�2��#�(�&±���oß���[2R�U�N�k�%- >!Z�1��dQ8�i����W~�:�>{9���$o����}�.m��؛���
�.L�5X�DN�y
���Q3�p�R����S
��G�r��I�JO'���fu����g~F���MM+Wg�;������0�u���
*��@�z��0$~��f�ad@����&��i��H�D��J7�vޕ	��Â��|f��^Qs )<6Ym� j��>dj�Ū͒�E��{����"Q3���U�D��Dᮊ�x4�l�	�C����D�m�zR�@x��rނ����ȳ׭�R&��H��$�����
ė�Dh�t��dj'�޶~U��M�tKx�1�[.�����8�]ň�/�R}1䏸�Ӑ�3X�;�.;�r_'�Bc�	� �� .֟�`����=��b0j�Ϳn�P@AA�(���2�(��a��s
�����a�F^���I��ߘ�UZПT�u뀇�gd�./��[�����P�W0�Jt�����3�2*����H7O1�h|�y;)�LآRK{���3��lEo��傓K`?�ΔL0rtL�_}%�)�՟c��&*'K����=�hTl�8^N�4D�mP` x�B�p�ԏ) {K���� ׽�Q�/+�	@�X8e��raZ'y�oz�����Q�pYF�"��2Y ׍��Q��E�ĭt�t棫� F�n��r>�<����oh� �?'���;��(�p� �N�ء�;>��A���o9S�����8O����V���%y]_~ou��Ж�F�-���\�2u��S�u{�_gM�aW�A;���a�_aY
�:f�Ὁ<��A�ܼP�.�E���$��0xB�\�!F�Io�|���BB���w;M̇���f�3 >5|�ʷ/2�������d[J���/[}V��҄��E�٢�dU��k먌/�U�����\8��N��9g�PY�[��d�������e4�s��V��;ğ�`�u����k{�F��R]é�'.���<�%�
��&'�`?+���0���'�v�꯼+�߉��ލ�;7��^u��Ppç�Ǯ����Bz7�p��o���l��8�6����oL���c�慏^���L� ���K��-a.��G؜g�=d;�p ���������1*�[)�=V��o��B��E����r�Y	�T����%�m�Z��#'3w�	���a����l���X���/ �i��rf�#j�齛�NL̖6�r�ϙY�O�#/��OS���`]Uʼ��>�߸����,\���H:}I��:���wϗ^)O��� �		na�Ma��f�'����=�r�~�a�P��pȏ�I����^�|��{?��C��g�nX
��G��V��J�~���*O�d�x�e��	�B��-��k�,���B��N$}3�ty����<�o�L���^}�aԳ��f����K�
*g�B�����]vԤ�"�$��i����٠䰺Hzo�ǅ��d��̤�^��ˤ���)��
���;�:�袮+���"	��rD���	�o�v�l�ӣ{Ox�f�6�O���&�=$xý�fQ�s2
-�nQ�BO��Y>��7	�����Mx�ט�kb׺I=��8�G�p{ʴ�}d9���a���m�6g'h�j_)�䱌�ӣ���z�+/�V�~��$��B���*ύ�8�����X<�f�6	�.�Dt��p��%ZeK�&���ńd��=�,���R��WM!��%7$���`�D���=���>\$��Q'2�9����U��oU*ć��gl�C:m18����}0g,����q~2��zUU��m�e�aʠN�EPG��B����Xn��"5Ö�F�i�����f�%YU�n�0��;���'�d�1�WY��̴�3l�a��c Lh�^7�k��lJ�PWy̥a�ΌH���>p�=��Х��y�iɡ `�����5�4R��,v���d��T�c�A9���FÂ��Z�!�z�2�r�'($���?���:_��ؼ�W��H���4�Zڈ���i�BO�<�Z�4�Kv��o�[�8���j$r*.hˉ­`���}�$s5q
UfZ����/�q5�zv9I))�LT�!v�k~�sO�u��{��w�`�4
9��ɞ��C��9!�Zv�lA��YPY�2�d������$IDE�\-��k��̒$�P�"y�c��쏆����r@��B�0��3�Pys�^�r��E��$	����I2SLϱX?ݑ'QMP��O��?�u�=z�@�V}��P�9��W:&�]}����kH��Js`���B��_d%ߑ�4��x�I�o2��;�e���3�iZZ�)G���S�I��j�Ft�xV�A�ȿ��[]}��{.��_8xLbhAp-6���^k^��N�kw��F�C�#�(Q /(�{/�� �옭�!�Cf����-�5R�8���5��j�+��L�?�:y��A`D��=��jϭ���Lz��'!�I����$q�f�Z㿻?�\~Xk���|�!�H>�- &�kK/�P����������"�r�>���41ݭ}�U-W���� k'�zz����&�O���t��Cd�Nðx�/���])⦛����6��_�ʒ�+�Y��"+�����G�^><�Q��8�J��jʃ��yIdv�O��yS�b7Z�8(��[�϶���?/y���W�|ӫ
�8:�.5J��Ea�m$(���:�pw��u�B���HMiH��H�j$U0bB����h�� %K�Ѣ�猶on]Z��D���d�UB�7�b#�Q]C���\{!�w������w��Ǭ��üZ)��F�c��U���Aȸ��w�9�L6��k�B���+�H՜۴�G�iS�
�\�p�n|�W��6'�d��Ds���gW�ُ�Ơ�F��K�D[$�?�1o�D�K��|y��mwnW=9����pT*70��g
�������}�L��n��%ȱS��j���e�]k��v؟�7��AC�I��ծ:r��Em����.`���;�Vg�g����3,��x�	X�:�p����<�m_P$\ߥ��Y�}�ï������Zc̏Y��:,�����ǬN��c-ࡈ��E�U�0�-����c�h-�N��]�(t�w����i�����S��%���S�F���I
�߶��-�G!���E<_���7}�@D^Z�捇Q�h���#ХK�Z�j}G��ʥ�x��?D-i�a�̯�0�˗H�7 ����|����k���JSOF9so��hY�5�* qm�'j�s=;��*�X�k��p���3
���!�_/(%WDZ1���
D2�kSS: AJ�����P/=�$�R���TB���I��~b{PK4R�V����1'T����/�A*�^2^���mÛ$u�o��^~���Ӎ]m�W�Ň��?����.�8��>"��r��� �9������1�0���#���V,V�q������D|�m��<@YB�O����g#a��l��<L���e�,	���xWoK1��Ǘ+����)Y������䯰�5�=�*rX�Hc2fy�,(O��-w�N�p�0���{���D�T�����O��̈́�eZ��/���'=��*������4U }1�x�@�6@�W2خi�-���5�_�s�:3 �]�ѮL����!����O΃�7JC���͑�r�YH9?������f�P�Ұ �]}5�I�L\����r�A>��o�rX9��e���d:Ba/Y�8�F�����%3ڋ�A�$4�X�E!&]���C�nJQ�9)&q�t�
�L��;A
�$E�xw����A�=w[�����R�����U�+�)��W��i�\߲O��0Xs�	W�^X�N$/�1V�����9��h��GĢr����M|m72݇.A�GrPQK��"�&'%ˎ�gm@vlg~�|Eo��	�bg
���������y�m��c w|��Aa_iN�������n|hE4�c�)�2�n��^<`�������)%*�1����P k�VW�����Œ/�VM����8�1$Y^+pm��ŋzdU�"�Q&�?��{�f�nS�Vq��P�ܒ�Ϟ�]�,.R�n��g7���ϱ�u�v�m�@��Ǧ�F�w�P+�m>":@Z���A��� @��謗hj���0�[G6�F�1on�s1f���]������`��X^� �h{��m�-U�M��MeH5?0c�!`���jf |yi~	Z��N!���������M���"XݠoXgη`���f�?� �F�P��7�Ip�p3���kQ���*��};լ���֟�=���nWn$�pq?��Π�L���zUw/3]�� bw��C���Dl�2��!Ռ3O�s������sJy?����p+�Os����Kxi[bB�5n� �bJ�^L#�R0�~�b��A���lI�1;8 �Lw�w�)Y�}�G�v �N�d��
�6]�)$�XSt����b��NKp�A���]��{fb�~��g���=�=�V�4-H9���i�+����^hG���U�z?��$�Y�����*Uzv�I*�Z�u�R�����*��PJ��$�,�F�le����!�p�k�B�K�?<�Xkh+��2�t�AA����a�&2;���`Kg�f� �G�yY�,�'���t���s����{.�jQU�sC��Ca`\��XTy�-D� ��e��y��ꊭc��9�(���ZW1�;<���!$C����*s
��p�����9�b#~8bL�������W���D�:�#%�t�� 	c�����i8�H��)/M��A1����j�!�ޥ}��YV��>�[Y1�O'TҲ�.�k��Z��V�����S�o�;M��|�'Y�%�� A�d6��(�<�^�]Ea�/��Q�&|@�i͚��"��a?,7���yK�#��aq{Ųv�-�[��=��84w/�IlΩ�]�g�.�*n{�՚�R#A[�v	��(����W���ir�h�Pe��)@��� 94ͱ�5��Fd�ͦĎ�{�[H�{�M��S�'X�a�ř�('�U�#^���R ��y~a=á�\O�U�7p�Vg��ُj�m�(�X̔��OU�l��peĒ�,��rp��m���T�G�7B� ��9��oNLZ?⑿����0d�1���cV���<�eO�=@��} �8�(ۋE��59� ���G��^|��u�\��C�3x
`8��vEX������
OB��D���Ği{xo]~U	S9� -�-{��f���:SW��D	�π���}%�z�j[�aP*2]�-zU_�sЩ��$��KGkBdՕ�[��r��u֖��|�|�꣣8 ޹!n,�+"��<w׺��\e�$;v
 �ȅ�R�r[K�C��s�з /��>$�uRI:�`�˟]�H˖d������K,�q<T�o���13�ö�N-�~�X@ZU*�tɗ���kM��b�����_巋�Ԅ`SL�O��G]�����.�p��.����V3;^b�M�e*��;���F\�XJY2�����s����`s}�,����O��RZ;��Q�����r�޻�����Ӿ�[�?0�ī�䠚s����d|0eb����Ƙ��@�b�9��GE)�A(��h�H	D�8rțjj��f�j^�D��`ƨ7��RKfC��}[��Ġ�H�ru�U��膊�X����'m����4�����h��,&�Z�+�>A�@��Ԅ
K���l-I��l���^]�ι�?z`ҨR�oN�ܞ���er�a�}�b^c�%�!fGe+`���f�'���}���u�K�<��7�r�z������rS=������rV��t�E獤M4�ۨrRRMT�������+q��T�}��8�(�b�/��w����R�C��81r���5��K"��݆� �A�;���p!̐*/�e��6@��#��:=�>�@@�B��m�{�T�)��x��ON7HR�|�*�=��d��ȸE�g�����]a^�%6�{�e��N=��_�S��8H:�t��ygR9&~��}�<�1ni�G��aը	U�|�D�W�6�2s�IȺ�g���y��L��f����[��_����F7�A.=�7��m��|#�I�L�_r���jc�(���J��ق��M���b��U��ǅe[x�1����N�?�C��ۚD���m`��V|K5G(3ԡh�b>|�gĸ��u��PY�'�iR4�W婗�ߡ?���Hek	��!�6����f���y"~����o'�
H�t�q�Os>�ʠ@P����R�f438���fB[JE8q�P%~��"�/l$Wb3A� ��r�����%���?mZ��QŬ5s�ƍ)���b���ы��[�s_i��@�K����T�H��:���1�\��emJop</DR���&�x��hM,o�f?B��+A"��
gi���}�������W s���Ѥ�w����tR�T�[��zX�Z����f�P�����(�.���a-۪�7d�5H�:��>���+��I�.1���2b/�SXҸ�2��}+�_;�Sw���X���G�����g�[7)��^O��sճOq%�)�5!~~�܄w�k�C�0����Y�E�w�(&�h	���z\��i�Ҿ�h�*�@������#���N���w�f��np�-��v�@b�5M\�,��#	�@D�Es����!��t��n�v�t���&��3�s�!~U���E�l���t�F�����gp�����w�9�g�`�J*5(��ņ0�O��G<�[�8�~�z.vq6P����B�GFݗ��J��3
��B{��8���A�����N�nX��F����ݤ$� S{�ީ�Lu�\��;��� X-D��r�ŧ��\�*E� �}���!��40'����g�d85��	��5���F%v�N���s�ذs�΀Y�	��ә����|�U՚\��ܒAK������;��B��1�]�yW�A���R���{��f��Fݭy��i
��2�;���>��IڷXx>!�*��	~�	޽�S�n��MY�KGa؝�
Ў��h#6�r��2�
�,�W�X�QfP��6�X�إ�,΋�[3���wX*{�("��v.n�F%�0t�m�AN})��7�G��˷�1�2�-���un8l��5��Q���ː��{o`W̒�����2��o%u$�b�\�>��s�Ҹ?��:^z�E�T�a%BZl�j�QvN�&	qz����@5��X���1�g���z^#���9e$>��f0�*��������R?�#3���@Thl�>�kI�Ң�e�!|�� �*�}W�KVT΀�����y��tm!B�u/�i�VC_t�LZ�9N�L���r��uPV#x =A:��Ο��U_@�JY,�
!�����u�I9}	W&�K.���+�}[pV�Tщ����ROD�جl�g���6���o�{���zq�Ѱ��3ȼw{�=t��br3�_���F_��
4q��}��	���=uk�(��o���!�t8tB���YP�m��fiS0�R����`^7P A��F3G��ճ{:x��Э�܄��L������Z�[;b���??�P���&B���8F�4�v��F=!u�ʈ?V�PUuB��f��
2�X��<��{�w���nt�vU��Ѥ��O:^ ��@����������)��N�5��O��^��i-K�8���J�`딵<��c�I�����v��߮9�WW½x�y�=H��S��������m��⭯V�����>nv�t��mv.���d=Q[�vH���9=߫��Y�k�ܬC��M���}��#Թ:����f��A��6o�#�%·���ݬQjM��C��&"��A��G�4ٌ��mc�h��2�����0�D������r.H��J+O�(?*/�?�ϵ�X˷�=��	��l.�ROˠE����:��IC���Ġ%e2S=ϵ���Q��r23�0���B���&�q����2�����-�MF�m����ԣc�Ffj����ϤL��G�+�4�v	��� ��[E9���t���:�r`����Q+��{ ��(�
#a�K}e;����F{�sY_���c�)��>�����eNY�A�� �6��2H>�R��*��>�[�!J0�Q�
����C��؆�{�F�M��zF}dI�L�Q�b�B�CG���uH��b��?h@ε�B�H���M0m#(�ζF�b>��*o�Rؕ4��vٰ��QS7��21mñ���?:(��,ڵr��_�U����H� '0`ti���`�M�Wlnb���,��IO	��i�T�F�rQbk����-�5.,f�i1J8�M?M�a�P�dy�iʦ�5RC����W�J��4��4�R���6���c� ?Q��$P͌�)�+��KQ�\�y�w���]p�-/t2$��?�j[�|'�����e.z:J�0��"�Lֽ��
2x����\T��0��{�Y��6=;dt�5�N���V�
1`��`<���ҭ=��|�E8!�T:AQD��+�>f�\��{ o��0p��U�Yߧ�T��U��ft}�F&I,��)�m���`�rjXc7�(�i� ./"zb���F����aМ=g��Z�N��,
cc�� ˼�@�g��d7��w{c	'p�\��V�ȮU�Vw��t�o�0��
�QQ9�AeY���<h_�랔�&�N�ȧ$%n&�N3WӰg8�WV����b��LW�dI��J ���ϋ_p�}���Ǿ��9�1?K��x9{m���#g6�b�_^T�roR�l ���|	�pxd`_M��y6w�̹Yp6\�.<S���D�
煳���Ԙk�]���y��MY}o>k�x��6&#t�ٙ,c���+��L��tǞ����D�����?~�֑�9���³�r�<ep2?����N�d)��4]-Q����0`,�a���B��C�h�P�r#X�"M�Ž�;����CQ}ӹ���|t�
Ap6���~�^a�7_��щ4�3�p�By��.3�5����"�`Mβ����x���P|����ݞuPYF�>����Ê���9�݃0���%���6��A4n��۾B ��>�Xmk$�s��k;�����v��#>W�tz{�%"��S�w�B�a{�܇P#��i��!���h*���v#��bΕ�cL�:�F�u{�^���?�-��~YR���#��E�����;�~X1�e�gB��+b�?�� �� ���k���d�ڮH�*� /"��b�'sܛ�#T��,.o��b��L��1�Aa��)�[g��m��-}��惷�� �ֶ49�L�	��R0ƂKu��2�,x���T�l�B��K�W1#�"b�u��1�C�4�����	2fFHb��m�q�&x@| ���͗]�'i�t��#퍗�x��+�iahk�x� �x�w7n1pG;~����������bk*jk�ߒ^�Pn#p�wA�Ea�$�������Y�ėa?�p-�a<ѶՓ�d�M������S�[/7��r�k�a�A�Z�{S�ٙ�|�+'<��S���m���E���/��#s<�b�����hv���s������vͫQ��ݱ�����Bֵ2����~!�ԧNV��|�!,�fO�L�!}�L�`R�ܐh)��#5F>.��%
0��n�y.�pUJ�%�q��@��:��y��<��i�����9@w5
R�HK��\��1�S������FOX����8���M��^+)ݵ��2ܬcks�L^��es�u�HBT���(��E1�����&��Y�Ǵ�H���;Q(93�i|.f�� =����8��z�g�	�T��1uJw9�_d���봜&�`�� N[z����l�M{��n61��R��X$�S�a������o$��>Il٤]a7��{���-z�g��)\_Mb�,`�E��0F���GWM%���e�_��X
�E��t�~V*JC4H�S���( �%�;���y�k�9�}Ҵd+��;�2�U%Μ�8��_{*������-vg�a�4�2~_&g[rRۢ��� � �	�=�3z�[��%�q�Q�REz�l�!���η˴�J��U7=D�W)qF�7��6�ԣj 5Kw6�c�e��k��F�)k�MO)1Zp<O~a���-��-��J�=��V�t��ν@����$���De/B*>�u^-}��xh�����(�wO@����k������+���7�\mt��Q��Y�%3h����燒���L��@97��5�J��Y@�A��Wq�b��v�Q4X%�*K1�ƿt�WA�2��N!d����w���S��F%�yE�Fv��H9�z[���3�0�8X�r�H\ \T�G��U+���j�����d�����H��r�����u2Z��/�T�h'�_�+n�)��'Kl��pE��Ll��Կ1{��)��#́���<r���2�n�C;N��"fTԉ�]�5[��b#�@���o�pV�u�6u+~!������9ܭy����-�"�L
j���ϡ�Nܘ?��0�=K^��wWU3��� �ڗb5��Y%,����!9��a�Zٳ�L���n��0��O�0�m]��><�����,�Y��j����\�i�C髏�i�EC�(��s���B,��Y�KHuS�]%��]���s����:*�ՠ�Q'f6T_�5uM�P��H1b�p%����dY��E3�c3�m ɫ���C��f*D�X:���m 27Q�ő\�H��󁇁���Ƌ���y�+1���9������[�b	A���t����-�Ě��t���߽�~o-���D&$Lͥ|R0��̛}��F��hr��+S4�]��Φ��c�&x���Rl28�s�K6�i�AlёVl`,��Ń�{��לu�B
�Gɋ����&�]��As� -�F��*%��j�f��Ae�P5`��R�C��������7,d	p ��$�sJ$Ҷ��W����3�p/=�>�-lP�]�5���.�G6�6�R� ���?R��]��;��j�Qt�OĹ�+X�P�-��85k/��DJL���D);m�͢6��T����&g��`c�����-58�Yb�EqE�~�冖��*�x��v˱k�(���N���ދ�ә���a��k��OeU*c�]w�kN�6]��A����`�fh�:J�i���p�� ���o�kLU�Q<���|���h1�p��Ol2��-,�Ty/�k$CB>��L�C��%�\�����pQ��2���K�A�8s��ҁ��|��A?7 �J���-j�Sx$A�Vb�n�Ӛ�Z^��
�*!~��{��L�~�ϊ�?�,������\�u�v.�)�O����c����zr�&e4�L���<�G�����m7"�R��� ^r����㉴5�x��J���:�,*�D��%�R"9��)8��L�e�t'rk#��p-���f�W���*��	��/ O��XOc����T@G��hޮM��q:�io�e�����	Gk����Z��/�n�b�V��BzI��>1�ޠ���Dד�3"�ٟ�f��jrr<����������Nq�1�D급\x�Hw{뺙/�>%��Ϊ��^�fQ9z3�C
�e��=��F��PG˽�Q���h��v접��jW��2��:)׾�=�x �w�^�ڟ�.�������\$�K�4�6���;�Q�|�ݾ�>[m�}�}
k�'�u�qU����F�y�UƒN;����ҭHې�������P�۰��v�/��{p�xǬ=mr�呖�L�[uk'�_�����h�j餸�w�� ����H�11��:7��l��?����|��!\6���ֳ���w4��t^߇��������]�?��}�_ ���-��˦1���,�U�����)��K�t."M�[��K`�A�AL2�ٖ3��&%�r+4@�2�1X;�؇ �����J�g	w)k���V��*�����ϩ>���W����a��gpƹ��M�?�G<Q�L](ܧ� �I�Ə���2�C�lk"=K!L����2l/��}�] � v7����=����KV�J�A��5���&!3��:�l�$w�?)���V�c�#չ�ٶq�\��ne�. �=�|�ܴ/���� �6I��ݏ3+{b��H�s��jw*}Sϲ��P~�9������(
 ��c�g� ��1y��2/X^j��ԝ��~Ӕ�B>��KDɫɘf,0�n�x��S��*Z'1�!�	��\���☛����Ӽ�K���fA����h%#RM�ϭ�;������_,ռ�N8m������,_�p5/�5@�Y�[Tjja��<���#�d"�U�!��:�L���T,.��q�*�Z��1��h,57Ħ����	��⩂f:�fL�* (�����1����P�]��)q�,�qeP�Ɵ�����!=�)����/	P,��,���mٚ�~s}w���#9����kcc��S��]f����n��|o�gr�[���̚��"��H���J�:��x��_du!�ɋ�z��Ŕ����)�$��v���Ts�΋�BC!ԬyH�v2�:�tw|�ג��'���y�!����_�yF����w��_��"u�������x�К6X�d�q���)�XtO��_�x����͑N�ؔ�H<FN}��6꥝���~D���nkL.����q(�>��E6����Y�\g7k�1v52���_5�dC�I�Se�x<�X֯��>j�_�{O��+� ��p����TZ�PDtnI�s��l�7�<��kA���/C4�j��UԎ/�� �<�6|�lVB����#�1-Ur��#�jB��cz��G�k��̿A)?U�|*L�kM�B��s��s�b��+��8Ax�VH��+#�&�Ĺ��������R�I3;:-�BPcs���L�q&�8h�փ��щ��V.ο�?���䱐�-I5�d�^㵹%�17���OB{ߡ�@��{���-W��nF:8���WUMn^�'J�U�Y��af�8����O�D2�W@����_��4f5bǵ����Q�;�[=�Cu�p.R��UbK�2�e�i:�4%��^����Ǌ�n4�F�3M-Zڇj�gMx�іp��Y�P/���C���8H�K)����=�{7�S9�<i95~�	�<����k��X��<vr�2����:���zg6A>-��)�/�k�Z�?�����	5�6�\����S2�'��2}}�4���k��23AעL1&�YΩz�}w��F>�$ǌ���m���5�;�$J�䰄z�!Д�织'�� ��� NH����s���Q$�O�߱B����{_(�B�E��MyV������
S�6G�|0��ఓ�e4C��� �TT��$�m4"�����
�^i�E�њ�YM#���;R��F�~I=ܙ[.�0@=�� ���[}"��i��x&�ݡ8�Vo�g>2��s9�\ޮ6�'?� E��ז����RN�c���P�
��~��1�}	��~���'i`m��t��sֽ���Uģ��r)q��ک/q�V�x_�0n~�h	���g��x)�����]v��y�\5G�;��8���_b���fh�4�䘢�����+�hθ��?��b��q8~�}���7�!1�З�)<LiNr̭y�6�I�Ve��!��_r���v�1����v"����,x"��@�!D�? �g+�#�T�B�[�z}��C���w���{S*/���7E�!v��ϴES3G?��U�����;2i�7��G%�0$��3ĝ��p8�!��l��#�Q�LB c��	Bl;�dPdY��ө&���Q���2��*9dT�.�v��9�0�	��?�g�JPma�W����QXDG�m1���?ԏ�rON��� ����k�W���I���[^c�,�l���[W:� �#H�kL���]4�Ƶ/�Q�Ƨh�J^o�_{0�o/���"��7�}A��t���"��[g�3��S:(|�����h��fcn��oOI &ڹ�g�d���7����Ad���&�#0���~�{Mb��&�+g/C��	̬Rv�M7�����^8RyÌ�~��"E,��!�u	T(U<�N��T�����T���Tc<��OU�+�E�<6�fdEƘQG��铖�㐐D�^���h�c�6�P�8���"�4N4�1�m^��/�)d�>I�[g4�x�kŕTL����3A�f�;��.��J�/�T!QƁ��)C��'RP�;b�f�D"�	����O1B>lX`ts-�`�)0�ڇ�6������"V�� o�Y�'����$n.ĕLh�����k8u/�) ;�o�k8F���w�,+���_���[Q{�G3L ��ZA�����I���di2K�+�2�k��cPJo�1�q��D(���9q#ba}L�2n=�Ŗ�r|����|�*+��p����^m�@>���ƶsQ��B���Hਖ�]�W�6�KE�#��o��֍�	Z��F������C�JC���aY��ӧ�Ņ����Լ��y���J�����Iye��҅hL��/���B�����g�Q6���Z2����!t��qY������Mۻ1��+���= �<��<#��b4 �-	An'�ceϥ�oƳ�y���&~_�a͋�'#l�Ub��a���c�"q�����_�>�cά����4���z��Ԍu�؏E&����cu:Ђ�	����x�F܌��}
t��;��>+������{N�遰�Sy�"~�h�旍 ���[��'�&K{���O�N�<����̨J�m���'n�Y�"6w���d��7�v�$q;�%�a���C�� �x��9�hm���I�p|@'2��U��/�W'��D��  gT�|X��hJ��Ý���h?b?9���?c��^���Ճ��;oɕ7FnT\_Ym4�56��"���la!]����~R��PD^h>�9�c���rZ��f�T��|)��$U�Ǎd˹�]���kݙ�2��*]�Zu띷���LB@l1X�<��B_"�C�a�Ez�'�0������ ��T_�[��Y*be�"�)��@6����;��3��\�O�\���öN����y! 	�1n�����)mgq�o&$vX���<�jL���p!��oyoU�х��qZ��H�&!�׷�o�G�*
�����~��:��M8��#4�h��U+�,��\�/k�"h���� � �Vz^
������~yøj�N�����,��w�1�悁O|p�&�	��
V�%}��M.�,�,;l�PekW��1���0r��NŃ���0�3��C1��U��'r�L9 ��	��� ��)3�Y{��R��'���6�V؋��r������F5~?���ah|��:�t��t����B�\�A7&U_�V*�<)1$xi[�}��IV�	ukvTGM�e��Sف2T؂�����S�������> �/Qt ��^� �!A�y��Hk_c��.E�M�%��x�L���l�\��p7��G����bD��W�g4Ɏ��OU�ߵb7�*��G�P8{���UY���F��#�Yύ��к����@.�bd��A���d����UΧ��~҄�yD5�%@���!���&N����<ґ��c�w�8�M��Ɩ������)�f�	��#p�2(
F��q����nM���,�A�fBW^O-ܓ����ݶܖ�������D8��ѷ��Ʊӓ�3�6o��|�+(tJ��&�⾀�#!�w�H�?~`�#2�сJ��0�q�v��	^Q@>c��[���US���a2
�*��=`P#U�F�8�)�F(��3��@��Z|�������8����:���lT���h�A�o��e�i�̝���i?����CUH�y% �-���\��)�2�R�W���c>�A��`��m���T	����Y����Rك&���3ǂ������@m�lvT|�s4<����.
��@�J$�qv��NL>$<��l��E���O��8n(�[l���r�}u��>r�)��˸�TA��F�6�A ˜�a�u���rR�Y�Gޕ؈-WE�@7���|���kc�۳ot���{	�ʳ݇����3������#t%�w�Н�'���*�LRik۷�YH�po;ĵ�	��|��
ߖ���[�&��7Î9zu�_��d~�Pc8�L�{	�F�h�U�_�!���Z4��.L���:�u�s�,��0S���υ�/t�I"�@���lx��5�>B��h���ʭ���G���-�xO<��]/0�7��[��i�tEvh����W6��z�Z����}0�Ĝ>��W.6���4��5�do�F06~��W=�5�]�kZS�2�\��9�ʤ�G��.v��?�`?�2�/�-u���:(~$�"�Q����B����a/p ����RŴy������1�X�F@
;��Z`�I�t��$�z���Q��;Kf��]�W��Zv���B��:�<�L��9(?$���)bz`NX��ĺ�G��Y��L��6Hم)@Fg�-H�`�k�QOX{I�(�y��vSх�_Jq��;��q�KF�Tΰ��.ݝvZ%���Z�b>�>T+cs��U}0��>tUE�9E4}�Bަ� ���pJ��}�C30�K7q}��������MZW��ܾUң)J�C��O�%��,��+ K�
����RG���tXбM1��֢_:q��ݓèlU�BNG�HK �Uiʇ�@�8p<q,m�䚛��0-� ���m���/�z���ϝ�?���s�s�_����a�ԇ'/1�<;�j����8*4v�7�%�j �00w9�tک��#3�Ϟ\:fױ]�Lr4O#.-rҁ<2*`��ª q��}�x��÷^�#Β|�ǅ������k�80�tW����lN�qᨔ������l�[3�k��l��-��x�X��R��L�13ɱ3ݰN�(F�sc0R:b!�SJ�7?PD06�,K!m���Sd��o.N�,�,��+���1)/�G	J딼q�&���+�)��i�jC����D6{�E����v���O.�-U�P��;���t��n�zm�(SY淋� %�N�=,��tH#%m����:�+�(��)��U����T�I��;��H*�M���$%OP�dV�.ǧ�C2;�x�}AI~�µ߯���.#� ux$����N�S��I�:��X���(o�PT2�܌w�E56݈>���E��z�e$�=�8Ɩ��:�݄%;�/�s~%�C���%-Ǥ�嫿1��Ӳ�U֕�U耨;�Ke���j��\�eOi�:�p��z���B� �2=�4�- �촬Ň��HQ��Q�78�S-V�uN,o���}12Z���,������I��-`S7Q�����][�z%,F��D���.&���i��W�|���+�w��$��_�U��&R��X�,�ĵ!���g��J"c"��u���ͻ	L�9RCR鲹o�0��xv��z�x&O�1-<h��g{&��M�g���,?a鍪�r���E��8r�VG������5V��d�Ϟ�}�y�5�$Ʋ���_��L�Q(@y5U�yF��kZ�eH7��ɴ[�Ƅ���^t���tqy`��5J�?�A'�@S(��s���`n��.\����8'�59��eɮk�q��~x��*��J��	wJqu��ק��w_m��z�n��Ie�:�8����}Z�i�nh_U��:����0���2�,]/Y�y����l�B��6�T�ʡy������j��~�OyT�E��/��ldgnyz�(��Ao�7����^�W	q���Ų03yB�
H$�Yy�ּ�v9�ϽZ���<6Ӽ�QG�K�Ƌ���O�w�|o ��MDiJ)i����8�lr���5���w6<�tg�6ki�=w."�J5y�|BT��b�A��K
Q��{g�O����)S��fO��wٗ�l��7:�)�/�r���,��x^�+ZZ�t������]�|���~�&s�M��ޒ6sh���|�Tr�
��L��r���C�11��"�%k�3Fg^��~���^�вfw�����ª ��R+�Yr�*��#���@�Q�e�����/�{�D<� �bYz�T =���g4��g)�R8�j���0Ե��m���nP�[,������Vh�(�r�R�4��0���Oy��q�J9* ���x�B��|h/)_������'��:�k�S���oDZ���6O}U8�*;���U���-����Q桐��i�7��u�-�2v�el�ru��ÑAU�-�K�-���6�W�ӫdi��)e�Կ8&g�⣕ʼ�9��EX/�&�9#G���SS�1�)%~K_��6fp�0<���/TH��64������jRÑ�@!_��L����$�����ދkc=�Hn�c��ʽ��q,\�m$�=��bk֫�}����3$0Rx&Y|�T��'?d�������,�*5���*bH-acw�2F��]�����-�C~Am7��p�Y&P'�!8����^�l��J���B�n���NV�n��Lv^P�c-��o�!�-ί��1bgf{�̽��{4Kx<�og!�� ����d ��~���lr����鱦���� blP�E�
]@e�5� +�t0�Y^�a����)�����_�l�i��.�HH6 �޼CC6Z%c����[��̞�DxC�,8��!?&��k¾�}�7wό��������7w~�z��_����Ab��^���%��=�W�D5h���ˬ��5��2h��ӭ��1�}����o��{$1��=��_�ai��Q�2��1TLA����VIxh�孑�Tք�1���<�gҿ`�L�f���5�]�:���m���\sC"5�׉�x,kds�a�~ 6`jx>��E���t�eqC����.�!��>�֘��7Ɋ�w����O��pCe�������Y�� ���IM�6��FZ�x�z��p�s2k.���0+���V���,�&C �}�k:N�ZI�u�w���La��������tnC�ʒ��SȠ�i��gٶ��h�@�E���ԗ?�.��׷o/�Y��5v���g'�FE�@��$;p����r����~�����Ȩ|�Kʓ	HH�J�[�G'Q���c�R^8��K�,I `q��]��iΚ�x����1%��A���!H4�!o��K�O>���Ӌe���gc��t]Fps&��L��>�HIo�'��4�j��"Z<�Z�f�ڝ�!u+�	x�-ڛoK��%5�h���=W�qѡY�׺�AZ�'�Y�dhXh��1�+�n  mJ��8���3��ƛ>�v���όN��[h����g�b'U%P�`O���&7��T0�`ZѣJ�p���~�39u� /�NΩ���䣣��9q�uDߑ������]�&�8�4`��)�W�5���?�/&玒4�䏏�x��p��@��'��<E��w[�Z��rי�Z��_���.�����I�<B�5�
�_�Avuey����}n�D >L�J��~~͝��p(e,!Z-�Ot�-}�M�p<哨ؤ��-��|8�J/E�Dߒ�]�j�ea��1�m�]��|��@����](���!R\���7���<�M���B#�fj\�#��j"^�Wӄ1�p���AͽU�"�x�5����l�E踆�!��|�F����i�s��|��y�i�SZ^n�j&Y�n|���Int���F��:J����(|�A���pS"^�gg��c��1Ǒjt���,)~�xʱL[����0�4�{����Ioma7Z��춿���}�{�up�P����+C���JYlo[�b;MC3-��5�,�� <��%��'2��7D�b�0G��������:����ܸӾ�E����"�&	��$�m
��B���f0H��kO�~ˎ;��f�f�Q�BH�FڞF ⌲���1��)P�N���#՘�=���rf�\��yI��n���'�ڗ�_3��#��z�:�F��5-��"ga���Km�|)9���^�N�]�c�_c��6���s���L��N��^�U%�����T"�����J4�'�"d�#铲T��5�S�`�*O[q%ʕ���ɧڹw�4U�����Y�t'��X���rA����'r=�N푹A�5���!�~�_#ı[|hW����u�� R����1��Te��[�)����0����J���'E��շF"�;�2�a�4 �As��*)�D�Iq���Ň��R�JW"�}I�.j���)��0v*m�<hn^R��Ex�}�pJ����FL�f��I�ϸ��-Á���ZB��N
L)�>��
�t�H:N�W���6#��c*�o�!p�A��8��Q�#RkZ�N�j#��h�����if�vXw)6����ǧ��ϭ��8��j59�dK�E��ď��6��YT�R��Cf�S�p�Cb���Ҁi�
���Q�}�U��E-�?r��J� K|�b<ͥ�krp�i�s!>'�9u],٧R?:ٕ�9ϴ���R��$I$�R�.pb�m��
?��ǌy�Ѽ�6�8�C�A�鬁��}�m� u�jo�Z'0u�����xPQq"{ x�Sw�c[����u`����н^6u�s�/3E�?�8��|�C�vL���qXr�zՉ�0�'�2���1�)���7�LO�������Gb�}��ɨ�ެ�NTh���r�U����.�:��wsU��.�^>����T��ʺ$)._��d�Oo��0������s8����j!��w�#�����'��n�L����h	��D���"p�}_�릶�*�~GF/�
^��KF4 �sN��'BSO;s�����j�5�L�,��}� ���	�z����?N���r��N(�9�񔈳:J��F��柔��3����o�ңK�4��N���0U!V�GM��缸#��N�Uv����6��X��:�'��U͓��\9%�j����E8�sa�3���/�����ѢԤ_Z��-sw+0�d�SĈ(�`�{���+�o|�}�~]���'d9ϗ5�"�r�O��_�JK��p��#
-"]����KW,�Ö��,���ٍ�,t�)f	=Ƭ�T�Ɇ^��9�` ��5NH�E���i.4ή�X��r�]��<$c����C原TJ���ck��u�Q2�$sLd�U+��]�'H���x�#n(U�y}�A"���]Pj9��~�#�eD�v�� B�t�Za�8�A���~|�����=H���к�k���5� ����^3I۬�#%�Ikɭr{�润[.�N���z�w=��-�E؛ͱf����$]}Q	a��0���w��k��"�C��B�$��v�\~�Î_|Zra�^|�a�1¹#0��w:YZ��*�7u�5��`q)n��95��bؘ1@��)�V�`��fp���|2��sw�LxT�t�Nn���
y�xT���OXa��9�-Y�s�Z�2��}�ꎎ�P�Ѹ�%\O�%�2D�˃z��~ޟz�%ƞ�l��$�(�Ȩ�kq��&/��Fx|�D�nw�F:���_��������<�?�1�\a$>�3���� �g��=��X��b� jz{y�(=���w{�����ɪ5�*�v�A�YV:��ܸ�aW�]�=��6�Y]aYn�%!k	�����.�-�\�ArF>L�E����͵�#C?P^�(���,jv�c��[�t���^�y]Sc�;g�=�*5b��E%�yH�����=���F��`:��%m�g 7�,	��"0�?sf�Fu2�~H����q�S�D�"���,��eD��.+�&�x#���x�1�x�9E��2��㤿���D�-240]�MwVU�5�'��ӳ���ǵ���_�E��N��M[r!���H�Zj��������V!�M�CV}\��9�0�J�\#~���ٛ������2���p�~��4�J��;�lf#y�p��D-�t(�GSL"�6��Fr`�w^�pz�f��m�\�Hޫ�O�/�6M`�(��/˗7��1a0�k㔢��v�<3���h,�'S7��+
F��M9#��#�_�-#�F"!Z@G��ɺ���b���jq�/T�:�@:w՝���"�2�+�f��=�LmO�p��_�X]���` �n�	�N6��Z�Nzi#�n/ϜB��U��~ѓ H�T�ܒ�0&ٖ��F�����6=�pۋg7��'M��2��x/��oO���U *�n����XQ�I�(���rm����p=�7 'NC~\���ن&�������Nf�O!�����>B�׏�D���'A��<7�A����P���z��L�'�a����{�2��by�Y�d7xZHv��҃�h��9��qW4�SͫL>A1f��TI/�����4
(3�8�g�d���:�:2ľ'�m�.A�W�W���j��b�q&�Of�'bYЈu�AA��ra۟���������4�Z�&�4����~�Ԩ�׵�~`y�u�O~TvH$z�\A0���_�<���0m����������x VGwh<�1��H�ziZ�y����by�2�Aq�ЌoU�w��o�V���S��CXG��y4y��c^7���� ��Z�P_�栉j@x��{��u�ψˡ�r	Y�X�1
�d�&�"���|���p��a� ��r>)���m������͞�Y��_�fa<�CC]s�7�Os�C���i�k�s�L���y��h򟌲��"�X�xdO���B�N��l�����Iqg"~+HZ�'��A������ST�&�Pl�x"p�m@� :C{끁�bLc��e�󯜗2OM\T�=�(F�^Wߚ�2c���#���>�5P!q���"���Դ/�0�ɐ<EMl�o���d��}c��nh��3 �zZU}��B�/B���>u�\DE��QS�,��d��{[R�TR���[(���&�2���mms����B/�*[j�iXO<ѩ�n� O�|�#D�c�Wbv��m���T��b+0J�IbF�z1.����l������
5��y8.��@S8�g�>��c|(�cA�G�|Wx�!���Ƌ��Z8	�',��0k6�^�~2�V��?��D6R�nM��Em1^"�!���Ф��Ĥ"�ƃ��H���a��.r����HH�rԈ�M͋���l�8%o\�
G�D�� *�1���o�	¢;��J�5</��n'�0�O�Fb��tk\�,�{zNjH�G��Y���$o�nU5&0� D8�DN��i���T�u�B=��U��bgvՂ�qҼt����/��\r{|L��x��^�Vl8�~�.�~��K +�VeR��(�d˺�����Aa��W�v*`�K������~ؾ/qR @��n{]���P4�B�X�Lc#T�>^Q���c=���;�O��ő)_�~[sT��F������mbuǲ��*�TT终G�j'lp�O�w�[l�T9���y��?����6����BX���gq1���]B����r��̩��vվ
c��G�:�1��厽ξb����HI���Y��2͂��Y��X�Σg�;�R����R�2��Q�}r��T*M�=� �{<��賏�R��;�;@�2ؚno��þ{��[���AmA��	no�ܸ��j����?G�����W ���ۭ���qDF��K����z�=L��ک!5X�x�wm�ÿ!�׃JX����F�,�D"�}nT+�8:���=� 4R��Z�ɯ{2-�F�t}�Y����Գ�2�m^Q<�w����^�x�m����(��y�p�B2Н�@��+[C��2�?i�8����N��{������SH~��쩓>b�r9���Æ2 ��9;7;�t�YӀ27k6DQ��0�w*��K���ؑ�O��m���J�x&/؊��B����y�& ����(����'��3ӖS@b��U��s��D	İr�K� �@��v	�G}��x.���j�C=�?�jW�Sm�=Y�K��l2��ܻ
o4w8�Q��2nO/٣G#ȼ9���؎4�
���Sb7���������E����.*�38#�4�'Ґ��.�#�w�E�T�O2С���s]�Dѕ�!���Y���\�Lȓ����Ւlj��Cl1j��w\���fy{�ģm��!Ph��������X����=��u�)�g����x�U4wj;&�Vd�F������`Үt3)<�)�͞r��]����+�@M� �r�4������˅*�P����" �y������DTkj�0����}+�o���aG�<�uѰ�8-,��٠�~G����6b@.���)� � �� u��E\~���&eihOS�K����  ��$�Gf��{�&���Z}�ӄlm�<���L�a��*�PG��4����9vQ�hֈ�tV��B9K|�o�q!��q	��4��W�WUz� ��3��m����L�v�7� JV��#O*c�H���c�ܺw��NS���U��~+�+��}OQ�qs�+�� {a<#W0}Er�LG��E����}6�@K���I�=�F�U;?I�jG�rt�u�Ab�4��J�NA�w���/s���y8�o�%�D�z&^�|zWP��͖k#�Mʗ���ԃ�V�I�n<�l;��6����߆�B��mЍ��X6F�Ef�'_1wSu��c8�%�pM�I���~ l�Y����<�
�稘`��F�kz�'��3�9*�c�����H�2��[�K]Г�tƟ�贩�}*y3p�t��~���ĸY.p�\��~�nSr@;����&��8�<D��.4��Ih���"ףR�>�۞Խ1�)���~�άA�M\�%��D����4
���R�t�z�ړe�F��Z::j����eh�/ �����;�����@�����^	 ����<�C(?�;U�"�U0�d���΄?",(f퟽����C�Ih �~e}B/3��g_��eE\�G���_���ŧ�
�?Y.���cR���3m�UT�M�EOʙU��2ϣ~8MȬ?�<���Ď�P��;,��T���F�hy:���S9u��ۈz&���'bCL�?&��vh���m����x5UK��鱩7�{٬��"��H���Ո̴U��RM#_�2{H�MeV�>OJ�*3����D�%�����|IF^E�Ve{�x���3l��������2�k�i	َ�}W �_�j�`��au(�����ō�:Je爑>��>O�lEp gӲ�S�'����{�@A6�%�Q=x�M�z�?�[��,�����4�����+/<G���&��1&NE,�	-'ޏ ~���Ǥ��iDK����j���0NG$�E�!G��r�)C.ʬ�1C�r�,T!&�%®����'G�j�X�©��ys��ˡ�d/H۷�Z����t+�������r+ӨB������0��{��Ǘ�-Gj���2�-�ˎ�1&Z�u6D�����o�����FX�����d��2/Ǟ��g�n���]1� ���Tv~ew,W�k�1w4aV�\�`P��Ӄ�Щ�}�N���:a�0�Q�Or�s�H��Yk����U�Ղ��ɖ��D�w֤�r���Y/�P|�������fz�(MD�Z�5���5�G���N�������2���OѬ�i���¸�CY*��MI���y��t���ا-Ԣ]
e؝���Z�*�)/���f�\�0pH���1$݆/�7tU�ô.�66=o�/$9g<�&��
�	|"���L{V�9�  +���q'\s+�+TG����k+�4��43�ᾰtk�����������v�!�_�o\*����8���D��1���&,Y?��:wC�n[�U�����<�L<bȒ�vR����E��[L�5|���+�g�: ��r��Y|p�-�<؊v��'�L�u�$	��U��c�c��Q�$.�4�ǹx�����#���P�3��8.(��>�v:��jj�i;G-z�a�dX��AF,<��� #\ ���p9������C�� h���)�T$��u}&��GSSra���g��ͼ��z�_�b�����VR[�����n�8������Q��r�)�s(w`f���[��ݺ{��B�]p֘9A3�@��I�'�$�,���"=��k�����.�f`��� ���~��-Q�\h�����pD�'^����2�{E����F�	i���J3fҾ�m;�9��q<����4Wu���/5]Y�bĈV��m��K`�_�2��V�B�v��L�t
��GqI��P㳫L�a�wg���;�r�~�m8mã�$��@�z���.*����1g5��a-����&������w����r��a޵���l�:;�׾�{^lJvI�1(˻&���m����߱<�����m�K�Zb��m��LU@7�5���Ҥ'���8�������������0�ۗue��
���L?���I���C�r ����
C5�^1[\�����X��DY���U8l��)�(+�5Vm�s��Ϭ�bd�JSa!��X�rV��+��i(]oţ�� WjG�w�4�#���k$���tEY�����>����SIʈ�����=,K��/I� ���3�AjU�X0n���=x�G+=���8���<~䃈�
�>�[�g�2�[0�>K&V�W]?�"i��eY�O�$p��kw����:D�L1;�0�3+�FKj0�ߒL�E�~�)�Cz��(��l��i���h{1�#���	~�7³���y��D��v%��`�s9n\û� �Aߜ@,ɋ�}��CSV��j�V��P]�A��H $'�]���'+�߱��������%�fn�"xx�q�u�:�N4a�w� ߽�Lp�Wv4��0��� ACޕi�����AǩxP�9S��u��C�l�u۹n�>�W童\�Fw�p>�P�>$���f!�-z0�xLt�eDyGʘ,�P�,��i�A8!���]^ �}ֻ��Q��`���&����i��jC"B.g��b�����P�&e�Ê��^���@������n����}l�žb���]�]��lK�<��G��e\�?M���ɔ$� ��Ra�~�]�J�Le<�GM� K��Þ����'�6�R��iA|����/6s���/���%'Ql̪-�ٯ|-��;5�����Ha	I@��0�$���S�:�L�m�5��g;N�z�Gt��
a�����4�~��0w��=�[�e/�$�g
�����־[���v/g�Y ���RTvQm�c\�#��'P؇���Q�(X*��
p�4��6���z�-L��#au���5G�+�U���~(y.���4"QQ���kAV':�p��e�i`�̌u��=��Y�D�����0u8(���&cf#QT�<��2�<�C�-&lF�E��wo����]Pޣ�y��6~��l�B�;��?����%mVZ��Ѥ���S��-,��5�$b��?w�k��F&;-r���O֗���T:O��%_m���<"Z����LS���I<���խpמ����c�L�$	�;�}�U�=S^�w]D�|��4��X��ϝ�>��D��f���z餃�w���!��WMO��D(s&e���z��(\buC��LɋFw,{��%���B��|��9�>��V�&x��
DI,4���6��jU$��Q3b^6lS�_Sp�ш]<	�&X���6B���,�xPz�̳��A�{E-����#�-����ZD�$.�`ǆ$vk���Mlst���YG�ǧT�YU{^ȣ��n�Aշ�v��2 ]#ؖ�]�Z�'-*�<�+�5"IO��3��	�U̨t�!���v$�B�]\@��ͬ��Z��"T"���T�
�F1f��!�Wt��6&E:�,Y��+֓�4>�� 	^�ङ��/u��wf	��[��E/���K�&1�MO��mJ��B.��h�=o%�'"MK����o���u��[����r�Q-����c��D��-��X(�U~/=�_%�՞�vF0Z���T�b�	�ݱx2e�j��p��'בy*{�����1� �%{`m���G��|�и��.z�ޥQԭ��io��'�rz�SȐ�d��2���F�*uK��@�
�q�Nsp�M�i�(��:CM4&'���	$p�on{b�ߥ��a(��3�'�\W&l3��h6��:n~Kr��5��?%_p�o��/��fK
1�
��$6��4��>�G�.��	zH>�P�!����G8��r�. �q<(�_���8|Db!�*F�Z��s×@��P�Sr)t*�a�b�%�X���A�s����L`q+Ɇ��x����?���g͸6:=�Z�õ��ʷ��p,{7��9�ݖC�Z�� �ɥ=�q�~;:��E�N';�|��K�2N,��g��_��r.f�B^��S�Q���y������)�{���u"z�1K-1�����e�<6Y�Z�|���@�"\3i��#&�Z���c�e3��K�x��f>ȧ���'�;��1�4��E��]��K�P����j3iW�����u�z2n!U8F��"�Q��/&a^���g��6
�-�~���(6�+U��#�.wz�)z�a�u�Y�[�Hc���e����������k�pn�T��z�<u�u����\?��j-C��D���mXI�ּdU�"f��zj���,*�!Ξ\ �<��x]���׋d�?j�Վn~ڋ�ѱ�c���.�ZKݖ��kk�UE+%�"�瓃�9����)<�q��>"�M�JĴkr��[�Z���iZ�~�d���T@i@�s,WA!�bVIg�����!�W�#�	�/?�m�3)!�a��|����"�Le�����V�>D�y�-�rio+�{�9BFٽ*;���\�W�"�P-��FL�g+�~D��_S�1�k�P�nwu����@���D��/��]�`_hs����0�L����fh���SF4�Dz�����pa�����.`q9�r&��q����ƥ�|=a��]2����J��*g���'����xŋ�x,�K��ۑJ�BRE'��lW��.n�17. �	 ���Z���m�s�I)��*��RԲ���D"�	$�w�r���{=�S�����*�~�l�g���rHK�eA��"@L�Ay�}}�NbS�S��Y*����r-_6�l��m�kK8{�K������8Rq0 d�d�;��WLF5�\6|�eq��Y�&Ҙ֫�W?hi1��CHz�k]���y����"P�#�ά}il��.�<�0EU�����ʁ�����zr�4�d������,Î�s�dtn�8 ����mk� �gh4n��
3O[Zc+)����&fm%�M�,�	#�X��]Ib�zR<F;g��/�e)�rB��_��D�h޸��xv~�nq��
b��j���2���l���*Z�����IY����"��5��|Z(�ןj��^���r�!�L&�5���V7�)�����Ɣ	t���7�E5�[�ӎ��F�@��.�%��ω	�`2%����[�kv�����"�j�h׋1E��<<n�����#���u�����*<�b��f�<!�}��4��/��Z(�����XӺ>d�E�Lp{.l����ߥ���si�Z�_��?���+b����l$��[��Sp��(���}����9
0w��u:b����47������v0,U��)�"	7���ȵ��>��Du�F	��b{��^��N?R�)F�?� w��������G1��pi���(Ng�L�%�?x���������𚥌P�~���^["4O+���:��V�6�FRq�d�:���(�u����&����+��Ӥ�8��M��W�L�r�d��5���M���ɵ�E���������2��Aw#~"������,��l0a<|����'Q�3�{e�m	E���e����^�\Ǚչ�9M~���]��\���K�|2k�.�63x����R+*N�)W�@!�Ey���cؗ�Xl�S�P~���8�U�d���(iԴ��s�,UU�!Ö́��
L2Φ8�"u�ܻg�W9X�qݵg�m�ŪR'@�����Z��w�{�U��u�?�("FK-�\�3�*�w9�� S��?�>
nb`�b, q-y��Y¾��^�?>����Y��n.��$�w6��:�����C
�V_�\�}�}z)s�P>���~���ꥏS�K���d���]t6T�/�kRIƱ1ڢ�Z�Z6�$ap�~+�bdae�g�$������h�r�'�?��Z�C�d�/�п��8��?�CeM��Ǐ~�ݎ�����e����y[��?I�yi^�->�@�r�=�ުh[�>��S��m^iw:ؑ}tuJ����|��WIB~�O/ ��edbS��z��0�������YŷD��<J~��,2꫾'.��ă^W�a�,<x�Y�3Ŵ2:��g��jD�x&�::��b��$tVU8�3�'��x.��U]z�cOi+����.^`��lf�@��Uxg��Zi?���r��DN�&V�_��v4~���5���B���i"�5˅����yo�z^U9�U/�2ޯ�g~ ����̂�Ko�(��d���^�)|��!�ey�˒�[Oz��[��s��qC]MhH��<p��
��u����o�:R��ҥ��*,��L����,Q�ŷt��� p����s��S�����wVGENP
��K��F�F�x��Ȍ��+�̉fl�Ө�.1���[]O*�}�p�ܬ�1��_�-�^�f�����|:эA�Q��z�;��C��/й�l�^硟�Ёv�߈�6L�w��j�Qx�Y�3o�x/U���<rh����iݓ8���/,|���%Y�>ݼ�������W��U���(�6���q+X�{��`��w7"��w{G*�A�'�6i��G�;���B�1�z%�M�R�`q4��m������(Wg�c�V�/~@*�2{�Km�L�R��j$���~�};O�o��e��k�-�p�Z=�$V���z�j���?ٯ(��} �l�~�j��I�l�R�]A��L��ٓ����@�-(����փ�ï��a�4�ԋ��,���P�"�#�(l�C.A��`W��T/y�3��	�4�	�U��P���o#6ֱ�N���	�V��	��n�-^h
AM?_��!_�0@4���aD���$�qڬߡD˖��v�riر���2���k\�'������M�vW\X��h�� L����q��嚺.Ir��\���=��Á��H%�g��5]^(e�]�迂��i	;�@ε���R=��?�I���N��/FczT��/!f����,�	�aӭr���Y����3�����Ob%��K{�}�\��y��������#q��sJ���Ԋ`�X��A�+)�vW ,!�1�m$��z#`�n�{KG���m8�7=��άц�w�j�u�ӟ�����-���j����������L�ڌ��
�����s;qi��pց@{e�2�2��/q���ɏ�iԤ��a@vQSc��Y=2�|�pv�hZ0򸚉�ز-ݴ�'�����z���+����; rv�kŞD'B�������h�$�z#�BãfA�E���� �#u��%I[���$����Opkn5;R�P�i��_:�jE�U�>�+X�Wm1��մ�̠pA��}��s
��q��e?�褪q,f*� ��Oݥ�n 8��(��G���*v�����������Vꤋm�^q�����8�ŏqƞ����5�y�O�~-��p<����")\��q�.��ݹ[t3�m�� #>�%9���YW�@��a��M�	�����"B�$J�jx���`�V�S"+U�e�
�x� 5|��ln�ݥ�Z��/�����`�sc�A��P >]yݡ������pB��^�}��sn�)��Uq�;T�b$�ߠ�:�C`YsE\���aV�Q��7$��=����"�e�v1��-v)7���ŝ��(����xiu�����ٮ8!*��[�zn���]����{�<x����(��Bol­�m����&�x�Gx�x�m��|�a3���%�����
����0 l�\*/������cd�s@��<�yf�C�fFۖG,���@�*}����2��m6��
�w�O��ii��ٞ�7�~����G�<�]؍#�ػ��N������{�b����b�x"P�0a6�q�U�%LW'H����B��Y�/b���؎bMt5��tӤ����f��������q�?�W�䬘o߸%��A�y�#z������G�X�	��J*��Y�=��*%.Y��0��~SK$���!Ԉ���NՖ�QTZ
���M�_�+-��t%���NB�Z3���Nqp�! r4��@�̗������C��öl�c�fP9��28<�o��lm5�nNlMð}2�}�?ȹ���~�'���j��N	����	|�R̙�7O�X6R]<烠	.��sz�^4 �� @�3ҟ�*��)�$��=t�D�M�1=zr��-�&�Ǔޝ�&�jo��(S&�GX�h����m�7�q:3<g^7����X�a"aG۔�	�����\�l"q�2�?U[��kށ,��B�9�����J���z�Ym��͓�-�CיK���d�[ٵAz���b�q���hg���K������7z��L����Z�&jX������-^��.����z�[�{\����
	�CI�=&�Oe$�"�P�����E�w4�b�(�����*�[O�[P'�+�ln��\��b_������ �~�#�	��޸j!���;��ֹ���A>�GM3L;����W��wD�^؁~�h��\������m�����"=h˳�z=���y�������/z��̠��_2��,����b��~P�NXHDi�=d�'S)���3�HY�W_��mo{.��.L�C�����=-8Z����6G$�nP��8<�k:X�h����4a|�w���C�LN!�9S��)��U(�2��z_����B�"v;�r$��p�cBણ�؇��uHMD�J �X��WD�~=���WQ�ﯓ���M�}IY��Nͥ�%�|t�z���r9b�C:�&��%�O��Q=�m��og��vv�ҀDC�3AEσ��9A�����뷕�'3^�/7��I��ņ�^����ƾ3W��a��G!�	��jzm�>�''�6�c����XW���r]n�K��b_g�1ү��aݖ^W�y����O66��c�=i�q)����(ߙ[B�M��+�G��?�3�OSO,�{�y�
W����Oō��$�VZ��~�N,ԕ�j��waBx5�h!������*l�Z��X@v%�Z���5f�H���ܧ�$���6frڧ�+���u`��x�٢PSx��R��)��6� �4eF�ϵ���x!��Y�8�ܭ�A��Z�;�Æ�?�����@��n���� �C�1�a#My!;H�����]��2��4 /L,��
^: I>J.H�*Ӊ�}U�I�cx�m�.�5WRn��Ig��[6�!*�0L��%�$z7��g��䗒�����"S���C8���8��=z�5�;�q���/\�X�[g�m�U�-Ez_z>>�b �@��1����,ꅾ;/)��C�����LV�(?Xp�	�0���ַ�>hȩM���ּ߁8F�v�:�Y���� ���*�j�*�OWj��_�,��4��ѷ��ƦH������O]=3w%ƾ'���f^���g�'���1���#�Mu��'n�������J�2/#
Q�#��P��kq�������И	��Hн�z�&�{E`y�����B�_�ƻ1 �(\���ˇ��,�P���ۚ�p��x��I�x0�����g�{Zq������cxy4�f����kӻ��gŎ;��h�J���|�2aZ��j<2���Z��H
0�4�#��0�	��^�#��q�լ��s!A�_�o�'ld�����Po�Y�tf��*�������}���l˾h�C��خ�åoY@U&�}}Kg�/X��~i�\���9���ٜ �� y9GQ��}c+���O;���S*�Ce��(�ht�_�t�%��b˴�n+��_H�|�B��<��g˰�f��O#΁�{W�����g.#�y��̱��l\e����.��F3��-$Bs���Qťem�a@Խzs����Ǝ.���,j��C0,Yp�����#Ù?7�J2#g�J�7������U�nߌ��Ne���v��e,/�.�
�L����wބ�-�9�&ܜ��`~��-b�\���VA��9-&� #ĮqN��n+W*��#m�4���D�W���ǎ�i���N�gO�.jZ� _�����eU�@UT�$G�)��P��S���+�� j�c�|�]m��/�ȸ^4w2�����t}�\C^�x��$<��T�Q;���5�8����;+������k@pd�{��^Q�Lㅼ�GwLa �E���ݨ�.f���ar34�B���ȫgV�e�ȳxFgzb�OG�W�u�c�7�G����f#�u�^��>��E!�+���[�����O�$���(B9WwI�f]^��4'N5%G�����g�SG�*za#��!7���� �U`. 1�?�u+�2bб)��֛	k������WY/�3(�5V�1�=�y�K�=�C42��9�_h��>���M�;�,��"Z�L{P?��?���zK88��zl�8-3�d}�������X���V�������az�s`� "�2pj2��Q庑�e9-��)�R��67�>{�)�Ek�&>�`�Tr�<>`�7�X����4<Sr-�i���o�ϑ�e6�_�|�GoW��p��j2*$�L�ķ#�C��?�W�:!��f&����������l���Ѻ�McF�6LN ���6˵�$��T//�5�3+%���3�Ev��*��^Jm6��K=�(0�`pNI�����5.��ֈ{����G-�� ~L;_���)���,?rD�Jb�����x�'�V�U7ܛ� >(2+�"�ғ�rUP�0m��4�4�`�k���Y�q���OĬ�/��0M.a����.L�J��yL����خ���SO#_�(�zAʺS'xy0�8{�I����BC6X���jmcu#����=/Ge�qR,�lW�ٔ&Q��{��&X4g�'�e9Te1NiF(�9���l�Yj�W��v�rA�Ά"��3J���< �����N�ZH�6��s����oY#��,��uM��?�HW�g�jdzA�Y�Ng���F���Z��)p�,T��X��["��G�"ϽbՃg�J�pj����/�Jj7Z3Pz���A���h�X��=������²q�p�6�����|)J����JO�AUM�Ƣ��H݃��.���;x��?}3��N���pTx1i]�<�Y�Z�M����yD�K�����w*��X�͔٠Ő�?Ks��Q��IH������q-oC_��;6�/������H�'&|�ڦ?�J:�d�"���4G��1�� J���.�������ulaTh}����x=�
�Yf�}Z��v��q�Z+1%���/x�[]�-#�Ve�K�y(�Ơ�����A����uE�I幆Z&�P$>�?zDQ3�NeO�������#�h9Bb�s7IŨ$���iV�H����4���KGՄꯊ���q�_��4=�II_�9k�N�6yx�Be+���֎ �K'�?=.8�5d�+��h����JTe����bP?cP�J��3�9��x��L���&bq0H������?(�X��G�	:=�Һ�<7د&�f�z���&�������#k9�d���V]�߬�K��e�H���n�`�x�Cnm���N��FM���ka�ޜ��z�ͺA��5�.%*��E�ΐ����n��U��~_�A�e|�3��c���˶�\�_����9q��%�Eo�����?��!N�����2��tA���0���>�ᬇ����;�0�{�&s��\���[e.R��?��ư7����Y�kѨS�{��9���Z�Y�c2����;A����9QO�V1��9���!q)*��v�71�O4x83��Z[8$S�9�[�)���ꢄr.��*(����!���6ǯlaCE�,�k
��\I��U3�7U9����Ik�m��*	1DbuXv��܆T�W�D�����{��R�ϳ����ީ�`#MUT�ch`��e��&�	��%\�R�(�<��+��S�7�	��zԋ_�
�[cS�e�-M/	3NQ��S=�杌Ԉ��k��� ��fW@�?�O�L���5(�`2F�wϋ������-�Z�_?D�p-tg<<q]�$`�h���Kl����GD)�og�N9���OkΚ�'H>����S���1+5[�����+���-�O �1�Ǵ��>� û��m���_��&�C;"��x�P������2��36�������F��2�^4��%�.L�n�����9'W���w�Y�A(���$N@�Z[�Z��ł���T3N'�g��A4D���|��4���������%J
�(�O���E��ĸM�:C��]�r�ojrO�p�c���̮�D8�պWd�0h�O�H/�%�x/K��5p��dF�(
s׀ �Ʋm�����羮���l��kVᄽ����|�|��b2�T�P�����~a&�t��/����̫�I��A�c�9n�<���y�܀�o��\L*IۘU!E�N|�vj[�#�~���N �G!R���]��aJ׎��پ:T�h��=�~]&�LW��0е`�ln0F��of�R箦'p)��|������7����OX��s�.�ae���PiU�zty�ۑ�|��?��m.4o����u�.�����LY���$Fb;�,������kn+��|"��=l]��B'������k}i�����9��}��`����,84�FJ�7��ƅ�C��d~�#�vp����L^��ϥ/�`���j�C�=R� ����]��w̽?���a,\�7�Y�����L?ޠ�R���2QzD�nq9���L,wF� b��A�H��h��4�MZ�/ �}��
u��1[X{8�����<�������i}��U[�|_m�^���j��\y}������VnI閊���b�z�_�D��U<^�m�n��'ɜN�ђ�Y�0�N�BM
Ԍ�l�Ik,��q!� ݎl;VM���3���O�g�O�1��k�>Jn{3�P�g�9-�,"y�%>ϳ� 	�Ɛ@!�'�oA���i#���-���8'�x�]������-^w�t�lq�,w56nz{"�p�O�o@�ȣ}�~��Z�ʖ��F��ȉ2�P,t����$�gw<��_��z5���-��.bq��:ώ��������M�,�b��c�:m�pPA�?s��T�uw��+�����T���4;�y��Q�w��;���a�A�I�R���_Ϟ�߹�p<���o�]��S׈��v|��|L)x���4t���%%c���=��q�ӮB�Yo�_܇ �\����S$|�	8�8`��R��Np5�CQ�Z2O�Y����c�ݔD��w��^Swxx��*O�v�:���F�6�^�$�9aqP#�Z8��?OV�^%�D]}�"G.^u6�t��F'���w-�6�e�m��/�귦�d�YB��T�,�W�h�IT�+֞e���2ڥ�o?�ܕ�䤪�h�6q&��I3_s�6D�!8Z���e.E���-1��ȶ��7�E�u3�6�Y�i�<����y�ꋡ��P�(�6�j�/�/�v|�N៮��{�hV6y� �p1��&��Ԉ	�
�����q�I���8/�%E��Z�@����������cɀa;$|�����k$�Q[m{�酽K2���/����l7N:}�����v���d-(r>��jŠג�8�#q\�������e5��=FS.]�H=TH�3�����ErA�g�k�I�p2�9Fr�j��}8u0��!n��)�%4�c(!�:u!^��D?Q�w��l�5;�x+k�'��wAC��Ls����z^�EH$��O�ٶ�>'�(PyU�B�c�M?MaV�"|A��c���xo�V��S_���6*~�/C�Ͳ��+E,��o�S�|ɜ"Tٹ5M�Qm�|D�uZ8��~Q<��j
�D������_��k��1=�):���^)�K��|#Xe�c&*�B����4�,BZ�fקLHCcx9෫�"�	�	t��@>u���l���9^�ٯ�aYi�)��s҂�m�?���8�R�) ��^��[�|�sW֗�]����mRX�Ѐ�IQ���1��eC@JaL�p��šB���cWa��b�����S7����@rD�7ϛ:@'����p�0UǬ��T5o�}:k>��
�Oa�X�ѡ�-,(��`�u�ҵ���5���3��l�5m�4W)Z��/����RR6��twl�n�����U�� qT�-������N���8�.'٨�Y���gp�1c�c��7���e^�K����R���	��)�}m�����,z�nPn`\�ި�.�
�5��s#S��%Vk�%m�on*>(;s��bd�7���u8Fl��7��J�z#ƾ\�bp�wC� z��my^��Sx![g�k����ٙg$}A�|�V�=��=����w�7�b�ϩH��	�}ś΅���|�F3��|�.v�����(+�z����)���Qς�����={���g�����X��w"��B&�����LxL�wPȯ%6]�r��l4��D�=5eC��<u��s"�dp��#�-S3˩c�э{�����4_�0��,W��&S[S7yd���,5L����c��B^ں������M�Xv z�jd�^�¡�y5,���5� u^��Fq�O�!%C�����V���(�0 �}�+�g��|�Շ��=Y}�O[�1��_C�)���C��� U�d��K���vK�Y����u;7bo�i�b��/$|�%��肺�*.��ON���R�s�*�\��;������HWW�ć��0Hޝ^�r���A��YW�A��gk&�;=����󈘼�>�i$���©p[X������kh	��~�8?�8SH�C�r��o��uB,��;�AV�L����ҵB<��v�$��,P�U|l��1!#�?D��zV8a�$��q'f�aj����[�1����1��W�8�;�y^�<z��r�/d/g����bƳP%!�<i����
�&j9�T�����l
�ޛ�Te�
wz
P��܂��!�O����'���$\	��4Z�@�m�k �^+
yc�Z���R�b�����_��\��V�&s@�N��*�[�HDE�����~�90��}SKݮ�o�������U����pd�&����]��P�ޫ�u��oh��@��#f�����o2�i�3��VBE��rP��#��[��j�Cif���6��2���n_�U�^�e�a�!�HZI�*xݺ�ս֧1��5|֑�5 b`���.�ޞ/���f���#��/����?����)���0-D�������"��PaT�u/�=�Z�6~���x*��[�	?q[�Y��bΉ���h�(��y���a��`fF�s�BX���P'8������_�h:1����g����>{���ԍJ�[r�iI���h~�`��E7zӫ�A����=�(tY��lɕȡ�j�jV>�����cM-�b�P�F�^j<Mu?�K8�4���/����ގ��>�����7��s?(I�?���-�Y�Sw��� h6��ˍǚƇ��a�;m9���^�>�	�~X�=$��tX�G�2�)+�3�7r��� ������.����۸�L�r�����lzG?
�ʚ����P��˃[��>h��0����n� ���[��M�O5`�3^ ����y@���	�ֺ�WNuᰫ��,.�L��������#%�C��
lHv�${#�օu�Cق2ס�F�3�x�}��v_dT�1~A����B�k���+��k�A %,��<zL�=�;�
�Y�Q�o=�b�h!g��2��pJ��% ����w�|��Cq�ƙo[Ž����� z����S9��n ��� �X�#���C�=��^�0�?<4�\ �E