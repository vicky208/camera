��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:�Q�z�n2�H�U��θC��f����S����t�P[�VS�K.v�$\�58���>��
G�]u�y"�M7/�&��4ypW�H(�����L�pT%�;6�3P�^dow
1�g؁�6SP>/�����M�&PXuW\yf
0�w[�MT.[�,�
����#�@��қ!�aD��.�5Y�V�Y' ӄ�P�HEπ*M���s5�T� +�
�%��x%-.E��� [�wj�P���.��������Oݙb�ߵ�?yh,�ҽ:pH$�Zdo2���S �%��5�������b�W�(�]�k��v6hp0�d�*t
�oƪɾ��-w��S7(9��)-�)(J_�aPR�����c�������m���3G�vL�f���c��7�Zz�0��}�fQ��-���9�g'�T{{+1%Y����C?�w,���H�]ـ��0~���닸���H&�jZX i�ig���C�j>ۊ��d�_�����9tSO
�����_�L7��M�Y�l�5DC��v@Eٝt����,r���_\���/�hA��Z���T������Pvǯ�P��;���
%vx�>�%����q��<��	��\�i
,���]
'is�����s�����,���ڑK�	h߃>�A�!/�+��n|���,p� �?i*9C�@�6��(m�1��l���u��G��u]mDn�g��[Tuw�\{>@U�����SS��aջǓ�����Ňխ�Y��1$��R������Ǯ�Y	��:��-�����q�($�wvLX�Sѕ%���i���NC_�iP]K���)�K�OX*H0�G��I7�c{��<:�A������uF<C6���Ʌ�S8Qju%�W�=��o�2R���5(��'�K� z���='Kޤ p~u������tӾ�	=�/��f ��<9��,Zf2��>�z�.2���HhkW�#����*���ov�E���J�\HNT�3¦��N ��v���mEK�%����)��#�hg-�/��y�Nߤ�|�Ŏ�zj5Y6�cQ:K��&��ѐ��e�RHx�
h�n��Ⱥ�C\�O��ڟ�CR����e�?�;n,a��%���$r�r��݅���/�_��ړ���آ�(����\�l�F�$7������T+��g�L��+Y�@R�LM��{�b\G�]�͂��8[]-��}�9���|�8����}�D��M�;o��*���Ŕ�7\�ƒ����d p�	!T5�.���M��p�����PZBВk��?������3�(G>�M6xj-�;|�Ec�-������g�bg�+�o��{�׌W_6�76�'�9������F����^�)άx4�j�RpZ<�}�-��y���#|�S0�ȳ�
�^�EH-v��N!A���Hr��М-�W������k��o�*W@�k�]������eT�r2z�R*[����g��g#Z����)k��`�X�n�f�Z�z͂m�Y����ꨆ�f	uz&�y��Rˤ88o�/��p��@��>z�(9��)/�pA� �@MM�;�'���)����YrVi�X���K�wo������b��Qg���0�͙�t�� �g��,ٮ���@-�rEx�����
#���3�����cJ#� ���NVP��$�����8�+��LnI��G������g��o!>~�h�鎐E?5*z1[��W-���Z��_���eR�m�L�	d�bbQ��̿�VX|M`Ρ�)��%�a>�$���E#���.�ÊS��0 Wn?����v��9��s�c��l��z"��ʜ2��X�%i쏀7���@z��Z�¸q���BJy�n�� �r�G�DI��]:�%�NÅ�L��_yR��L�>cꈾ�<��*k����������]�q<�n��pU������RI�T?�~2mX���ŏ�����o�hi�b��K|�E�	ٕ�4Qm�`��I21ZA��'^�<:�L�I��S!��g�������w}4�C7nO��l�z��-Xm5ѕ�ԩ�;^b��Pzb�6�x?ʿ���
	$��ǋY5*W��`mRQ��n�C%y�������-R����ex!V��\��2�(F�Ah�8	K<��|� `p������Y�8$�΀&z �W��!#,V���W_}�L��1���>��O�܇s�iO0�8f��C�{�&/�
�|�`1I�Exg��Py�}Τ��l#�ԩwRM���l9N����fX��W<S�Y�'���ݪH9���;�߭$��{j<����w<�cKF�׎�y7lY4�g�n�s|Ʒ�T���� �X�it���]��#B�ND����ݛdڛ������
]C�M��uy�C2<˵���h��z�ׄ�7����|H/zh�޴�'(ܭ8CX#%���b3�LԦa
�1��*�Rl�lo�L�0ۊ�[)3�VT@��[��(+\\YQ���d!��
�ͧۜ����Rѭ��!��Y}�]��ww�<}$D}���tܧ�m��r�)h���gN>B@q�1Y�I� �N>x���=�Q��'��\mt7@�ŨWwU������.^��eĵ�
������~^�3�6�Ug�;薩�
Vߡ� !��+���V����HY�#D�g�zb������X����|#�)kW���M�xr/���z��X}�	�o�k�% &��'��
��c�wE��1`�昋u����1E�|9�9��'����ZX�3��-yS�,:_�o��r�m��f��;0�g� D��Ӆ���Q'O���{�4ڽQ�ui�";6�Z<��G���)@�ߦP[�H��2��e'[ź���}W��bƨ��#;P�"�s3�:_y�Fa�(����b�ۚ�Մn�������׍B)������
�
�h��W����"��=R�e�h�!�B��ݩB}��ȥ���P}2?"+����-Okf���4���\>ޕ!1n�����Y4Io2������`�i�"4�����]��@��Q^+1�#՗��e7m��yu%�o>����Ze�	�l�Nz��&ߞ�<lv�r���I�N�y��إ� ���=��)٨��	��� �7�����4��M9��9ͭ��aw�`�PH3�&+�8�p�v,��������~o@c���'��1۷��H���@ڟ��2[��42��ڦݖʿ5'���Yt�ny�w�63ނ{=���w�R�ʌ%��J��z��� F�j�����X��=����x�0�B�ea4��Y�|6�%i."q�i��z�Y`�a���4�����yT 0;���v�n#�.ׄ��nA���c?ר��ƾ&2��xi�R�:���6�<���P��>�4J�fu��9�3|C�|��.���+8�L[�[׌<|�8���;I�4٭��7�(ܰu�g�����	�y�R8�Z��Q7�;b�-��[��ra@��@O�D�o�	.�4+��1F<N��'�Ļ��шn��jb�����(�L�\2�Il�wTL ���PG��lԡ�]��N��l�ۏ�zc}��}9�&G䅷�`�D٤똂�X�լ�^=���&�a�l���Dm��C��}����(R1I\���}�r5�O�^�<��agZ0�M��³\�	3�I��(�.��`��Sxk�S���f&���g�H�A��@���I�f��� �2-��\��44� B�զ�Pጮ	.�<��8~}O�9�Zn-ŵ�)?BLZL�Q�Ƴ���n"�����JC ^{(�#')I���mo3�=�MM�]ӕb@��<"B��d�aҿ3
�e8c��xa�eFaT��Y�r8�cy�=G��ȕ�woAE�@k�����yA��"V�@qM,�� �U���y	Bj��[�5f/��� g�d��[`��㻙R̥j��۴��ft-ʏۇ𻀺��l��S���u�����W���Q��̍J��֥���8����Dnb�!��նl��9��h�^d%^K��V���{�& ��rS�=�E1��cT4~��V�l����˪D�x�nK�CSr?\)���&;�	�W8�_���7S����d\��~����5�"��� ��R[���U�t,h��&����<)�q�5'�&X'�r�I&�q�����跬�o��k}عv���Nא�C�x%��i�*O�m\���'��u���G�.��m瀪v�i'�/��G�v�%A�Fi���p ���)B$���^�nk�߰�C���C��"�7�op�=��o�ٕ��X�'�{gP�`:[tv�0���h�O��5�%���}՗~E�@1�2�ʵ��Z��NA��r������mQ��W����󶵟�@@ݘ#;��?�����P��(}����E9�G�����w�D�P�ɐ/9녑�xr�8��������0�k[�f���I0��Z��"7��F��ېt�.�!>��/qw^�l�Z�^�>���&J�W�
9^E����6A���lu�ܿ�_N/�и���;�곜�?6��^f���q_'"qF�fW�Ơ�b�c���۸&��:���Z2g����ER���q9�>���
Z��l�j</����C�	9�R��]�;.ɛ!ڼ*~��O�x�8�8�[�ȏy���K�SM������uw��n�`8���r�[�N�JV��=��=�8$h^�+V[L�x|!�`��͸�a�χ!;N꠰Wi+�J �8�bg�Mb��*~�¯4��,_��*t��-��a6ؕ�*�-�ܹ�S��^���O5'իN��<>�:J�]�~�mdd��*�}�N�0����K�U��j	�#�3�(���(�G�[�(�dÜ��M�;��Xe'C�����p�Ƙ۱�C��gPn�.J���ty�8b��/��k���('�r�Y��#�$uQ���r�N�`j>�����m����K�Ҙ����BH�Z��)�\'�;�ȝc���S���cpq(���;��닶D��o1F-ѡ��&�� O��\'Ȗ�č������\`,e��U�p���C{�c�qqf����龦=��/B��f=s��
I	��^���l��2="���ݗ���� �N��w��95k�^��_�_8�h���������xa�?K�!�I-�3צk��mG1&��"��
Ky�|��t�jߗZ�������y�?����� �.�P7n�����3�CYV
B��	��]��}�S����\�nJ�&�9~k���z��]���)�Nz[�[�����d"­Z��f�O5]��S�!�r|^a�񑡢��q� {8 �����^ _1$��Y[c������S�n�ݹ�E����
ޘ�\�N|L�������' �ۇB%X�٬����s]f�5ì� ���������
/����Q�����M�~�1kT�cy3��ո�q[�ٹ;�h9�OJ6h$g���2�.��ȷ��ʸ]\{����G�H?�p��<OY�_��G�u�z�!�e�@�p����mA�ѻK�4�����o���"j,5$�fBXn��9eΕ��	m�3���ǋx����^5�PK?=��5G�m�zv��n�=jL�����`{o����
-�*�'])��{�-�}�㭶��'����F;?����uN�Ël���P�_��1J�zǺ��`yN��'�'}�Əg��/z|�=I���h�a�v��EC���+�nޕ��ͺ&d1��:��k��Ia>�.柬��}�������Gb�{MHPmbVk�@��9��W��gTw2�n�b�s@�ԅ͗�����)�_E�$n�K�������q�L�e/pJ%63���!��0"ǿ�N<�ĀXvZRO�$�P���K�!�I�`cF�V���.{1�~^�w
`0�m�`1�S�X�|��,1j)��b�S�b�@H�w���<ֆ��V���;-q�U`�����+m¬�2�)���)9�[�TT��N�����ۈ��ŽG5���V�?���u[�!�]Yhۙ{`��CWT��م����'A�(u���G)k�@��!=biV.�����c�`�3����9��G�ʛ�m��(��%j��5hCS]��tʷ�*��������mǘ��:�ǻ�-QA���D�)T��n��u��ZH{�Hi��ᯍ�m�����-�YM�@��L�<td�Nv���D�b���}řg^�ՠ�n�N��\�2����m�*�zM�Q΄4-
���A��{�O�����O7DJ~H���=�Q�p��0��@���:m�Qx��3����_��ԅ���؛�sh^���j@%�.M�W+��-��9I:%t!MY����5��U,�K2zEe|M�(�q�R���[MN}�I��~��$���f�� `��7�T:{���Jy�ۀ���BK��b���4�'�.*d^q��7B�̙����m	Y=��(r�fjވgѣs�ݿ���SY����K0f�-Zg��ꩀ��&��!�`%M�d��ß��9�|�UNSr}���p[T���F`���'=�	0�� ��R�{�����w�"���΅鏄)�
�6��?7,@e��l㛬�I[�ϰK������t�}��9^���x[.K����@t���G��Y�U5!�eL��%��g[#�����Y�@�Ğ2�Z����Đ�͝���E���f��0�\�p��vԬ������O}8X��"q���g��ب7��W�R��\�k+��: .��ӚѶ�����Ț�P�z�;$���/\T1o��"zx?aP��hJHݸ���n#�%��)�@bGK���t���H��>Wߔ��.\�S�3��c.��<��]S�T�@����Е���8Jq6�`�|�ʁ��
�@�#F�G���;´��O?,��Z��oy��d�F�2��-!��XL�������ҊADӲt&K�k8aE)�[b�r�G��kg{�?��$I��h��A�z������F.�]B�^�6�gVA[�է*�����%��g�R���Q�O��ٰ*��L���8���@�d��]pS5���Tw0d��'�dCa8�y�}o��j����A6[���8Mǽ�5���>-A,ko�fJ7jk/9Mi�h����:i��&���dK�\]�S�B�o�V̒(#'x�M�����_8O��~�����K�hޅ�E�΁bvs�� ,��9����?z���'\J׃����!�74����Kg�V�ޱS��V+�}��	��}R��k��������h�1���'s��ʚ�
���;�[[��<+��t�Lzzc#�*��5D�cΐZa�O�n�_����F�	�fW�yp?zKJFyWX�/g1Q��I�sx���;�"	���5�!x�Zy)P��O�߇d�h����<��c�Gy�,Iv_��L�����7�������^��h_��Y�C��&��B�=SDאt [v��0��� $�\-����	��N��}���(D�Y�sPE��/�ԏw�ТF�J�-����j~MH��ʯ��~�c#�F�]$�M/��m��p=�$��oru�y��&���73�©Aʉ�>�y���5(t�94~]Z^�dQmd��,J2�'��\d��ဥ
�
HnaA-�������t����l��DgЬ7f�Y�Z �{� ���Y/�r����&i�"Y��P蘍Z[�}f�9�����cv�փ��F�g����F){���*md�;rT����s�K��	_vv�޻�f��P)�n�az�Bxo���������k �@ʓ#Qw�_*���?\!��`�������|�à���6S�3���S�Mp�1xK*sŐ��n�0"���4Հ&�(��a}۹x2Ĉ�q@ȿw�?i9^g�#;k��2����)�d�f��կ�����g���|��j"�����!_~�͂�ĝ��jj�c>������J"ܨ��ӵ���\���lWX'����f���͕		W�ޙ�X N"J��/�X�U���A3�L	�ܑHC���g��՚�����z�T}H��Ts}
�>DD݂v����ͣ�X�o�Xq�;�L��n����o���k2�������S1
V;[�b�Œ�Rn�4j4�W�L3�_����Vyg��8� ��Syp��Z�owbZ����X�Й���QP��7�>���vH�N]��gI%�-}�oD��`4�2HU��W��� bV�s�|��~�y�И48�*9��0���?#G=���<n���T'�E�{ckŚC�WI^��:u%W��U�MO�΃� Ȕ��3�Ҍ}*���)ǖM������t�XK+1���D���s
����3Iە��or�8�V�����V�mʠ �+tƅ���?Ҽ�$��D��Ga�q�#���5��L��3<i8,�7c)�M8�V�Ze�¥(Th!�깐-��J".�u)�D�s*��"��DBM�H�V�~�H`���V,=�cfC���j�����󂒋YK41�5���%���x�.�uhϲ���A��i���&k�0��gu1ύa)(�Sv���B^�(�:f��cO#ɝj�ഌ/�6'�LD�N�p���X)��
����}�[��-�X.z=7$��܃ �A��/���Z,'�S�w�M�w�����l��FH�^R&�zy�bN{ۆ�m��ІE����=�JHT��Xj8C� i{�l��;zT���/B�9#��Q�0�uR�$�)y�C>���v����S=�\���or��,��&�Ws��)Lq�kl0����N�('���CZ�a$��a#�3w.��a��MԀ�S�*�^|��}(���-h��Jm$Qͭ)x A-x�H�w�o(�K�\���FZ����,�S���W�[��7����>����u��w/�5���]PҎP������������m���������8=�Z�o�ׇZg PD�%K�]�-!Y�:"�љM}lP s�f��H���mߏ��r�|\A6�w�P۞�`�'����xeϼ�ˎlg�T^���#��x��Gm)��캘�, c�����v5\���6��%�w=�H�R�����s��9����o��=������9����ǐ�X����빲ҦjZT��Pe@�����?�G^"�}K����;�Đ7�L�WŪRp8c���@I'QL�X�ө��iE��/%炼��f���#��j�� *�!��̟�k�2 dM�)A<�9� �������3��й1���2"����v�=[��<�-=;�>��l�Y���4?(�|u�R ��Kg��5qӽ��R�W�&��ܔ�mY�����=�)62�{�l��FiZ����Vc"�^�px1�{��NNSF�!���$�D�˻���,9J%�p�� >02��ɦ�)cb(?o��`z�����N ��o�G�}�Bmb��2���X�w���*|�g�g���y���EF�Q�R�d^��.?���_/B���9"��� �0���)P�s�|H;�heH�xpTG�H 8��t�Ҽ��͒�gѪ;�ow,�{�v�Gl�� 2w����Y5�H�}K��)��Y�����+�;+���S_xH�/�}z_���qW��/�kOĎ�.���)%.�ua:}V��Wnt@�͉��"'ؚ+�-�\?��F6x�k�X�VS{l=D�5O��c�w�^�8�q9����[������ڦ�P�ln���y"�ƺx�
=��28W�j1>���'~Gm+�����!��dHg�����5B�C�]�����|^g������X7�I99���ذ��=V���>�׷˔�j�?G��BG*�Qs��F�+���H��1�]S��Я;~�SK�gK0.7��P�%�&�.]���	�Z`)-�4��S$��zL�pl����yT����WOS���K�� �n�? 8?�;��<}�6���� ��N�C��|��ť�ss�����}����N�ֵF��~1"}��q��Ts���@�;y��|b��[��\��p�7u�P�7��«*mMfQSA�+��n���.��q��y��AF����ehM�������ņ�X{�K��Tʼu�P&G�t��+#��Pl�Vȡ���;o�N;z3�	�t`�E��!��7�IɆ �� ����.ѢH�	k��u�(<�Y)��0� \n-s�I�����r�5���8�ɟ�7��[�zDCzhQ�]&/y��BO�;e�4���);@�!Iپ ��d/��%�"�8�MD�K)�Ԡ�1��l8S9�?�f���4@Yq�vr�y�y Á�OQ�g_h�%�ћ���}��O=
| �,'˻�H�ݿs<߬�[�?c"(�Aɯ��ի��I��a%ܰ��o%7d;�}q)[����F�H���G��-Sh8C�+e�أ���6%�`��rP1���VRV�����M|M\�2��ȶ"��WR)3랫&&1s�F�Ϭ�
�Q1�~+}?����|�L��5�uln�UހΆ�+�S�H� s��t��pS��Ƶ�i��)���Gg��+WX#D�����!�+�s,ŒBଛ�A-�٣��GeX*�[�āȮ��h��M�?��y�D��s�c�H���BG*9U7����]��V��A
ʊ࣒�Ր.5����z�K����û�*�UF���,ɭ �u�k!���L��҃]ꪁ}p�Ut����p	���n�qX � ��!{�����}���=ܪL�խ������B�[�rt�*j���@���LqB�����~�F�4+0T&��w� �ke%ˊ�D���\-8,{��,�i1Q�����8����3�ͻ���(���4���W)�4v���!���q*5�mB��Y�"5�@51�����"�/�{):�u��y(oЧ^�~�W�(Ŕ�
��_(���U�O6��b��Ϻ��d-�5 �,���@^B��n��翵�b-�f^٥ˡ��l]�C��:>-��5K�Tn͵�1*���K���-�!����b�u��	y��bY`D68&�n5�F��֚�;��3!�u�	K�W�	���;�W���(⪕�)1LO#��z��x'R缨�����2��2<�.2���$X���I�x�W;�DDFk g""|��i[m*OZ��@�I�	�vX 7G�z|F�[D9���|�z�J�%G`7�WǄ�8~�M��č�V�QŮ���q�eM9-�oM�����)\hf�� |#.�bh�y���pS<�8?���tG`��Ǒ�T}�0Fi�>��8��q^[�� $���B=�@��<��Pvk������:-!�6�_z�a�:a�GZ'#�;96��tGEjS� b�J�G��q-��z--��!Xs���q.g��C6�r4��4W�_�S��B�t���W��la�J��p�XPO�[Y�VoO�+���
S�Jh<<��T�G�>t3���K�'�� �z_nP�9?��X?������@�f[�AoT.�)@�u���`m��Hж��C���ǧ�'��N:�*b=����_�(�6��[�6��.��(f�:o5��C,�,>.� t�+ݶ{�H��u?�_�b��̵M�I;r�S�"��fN�yo٣�y�4Rϗe�\�Vg����%D�qpi�ʼ��y7$'W���ٵw;��oL����is}<��^���b\v.nK��,mME:$]��+6����v4H(�[�մz:�ph�9ou�j�
��Ѹac8�u0-�g�1��y٬�7]*�T��R1�deS]Vh=
���}�|��ϕu��(��@���lp<�O�(X���z�p#&�6R "�[��c>ǲ��	�XbH�M�M�Ft�7�!9v��Mǹ*��M�˸��xH�
h�P	毯��}��J��Kn�Fnh+���b����3S����^�w����H���D�\��/��x[�W�Q��i��	ô�#�����Unn�i�	��j0���V�g��TZ��/+>��34���5�K����/q2Up�ȭ[L�'��ƭ���� ~ދ���l]��Tj4�ٕ�ͷ��	_�î����z0E��7�\z-�1��OSp�Aր�ӽ�ׅ�H��g)�S���� Y�i�y_�9[��d�^�	���ڌb-�'���#B�t���1'^����	G��ɿ$U6���{C��_�lbr�	����5�'�h�e�R���n�A=��ʐ�NˏK?���5F`�5&��+�3��<�^�������C9ð{��kO䚑s�{��e,��Uv"]�hЦ��w����-q���F[�@1s�)p��Sq^�I�]b��(���w����ܔ�����`k�9��P~fQDl��4���
ݧ�����z�#�f'~� U�H�sOu��O#ïj�Ƴ�oY����֘s��=������O22cR�0��*���E�?2���y���tw�p�d�O%�W9��d�Ѿ��̍TtY��k��2������w��"�2���y�.��BVL㱐B�xὃW��1��o�iGi�C{���E�0���U�H�{��.1B�?��߶����{�*��E�6+�U}����'1پ<���˛Ç��+9!�b��/%�Z��ޅN�z���:xk�]r���ʾ�Jb5Q�rՆ�'�Q�n�m�B�D���������� :yB��U�����+}�39s�%�Z��{�"�B���r�Z"��L�� � �A���z| �;���z!�c����F�� ��<�XD�`փ�}k�Tv�8��y���:t<�Z?;E=�"^�IAqi3ʴ$26���cϵ��vL�c\_����[^�.D�O�5 e7��0��DY�@GO{�is�C�c<PF�LZ����V�mzQ�쯁���fC|���}�Xτ��	s㴂�MJ ��ڗ���Ęo�MFr��$l�\!��q�q�5Sg\�v~X�-D3�\�M^/��#�� �)AQbQ^���k�����E@������d�˝��}�@�.�^@��
�%���mw�G������ob3����)�;<8S�l�?f�Wc-�K�ʥ�D�t4$�N�q����+92�3RN��!"�ʹ���PJko���P�3�i���7�ʖc��v��.͓�_�J�Rl��#}�7=�������N����a�e�_Z�!h�J�ꂄ��x{8᜿���0�v�3/	�%�I�J}>$Ez^:�V����Z�Yd�J3�U��K�;;��3_�L冢� ���lO���?�:s`�u�5:�x[����H[��T؏]G
�L&�il��A�1&Y#c��~�kZ�j}�>V�<�ދ��3�`�����_�2�"���*�^u�<��w'�"|�����^"��~��uW�6 V-�:����^�w5��z'x&\�a�Q�3ˌ	\�cqy��ʼ����%�N��(ζVsK؃�����R��1e	��#S���L�3�Q���(R~<�xǐ袀+�f��;����S�s�kdQ`GZϠv@�f��^��q٘��9O��L�=:e��E;V�VU��K`�@eh�]�#��š9ސF��k�$��Q�/�#<���Q���M�����xj�Y���Yc�J�j����'rE�(�Ts,�cjEf�ei�?�`�hn���.3xx�ncݭF�I��������1�ni|j�q��㞊�N�f5b.Ӓ�-�@�Ȣpn���䳱.ˌ�2���`��5��n�Z'����ڙ��c̱����AJG�ƽvU����2=�߷��2f������o��/=����VXD=<8C���3�0ݺ	���X?qG��$�C2�ܸ�/a�կ�Ά���*]I���DI������qx&�P-����a�-ek�h�Ǯ��ܠ��8���4�YUR��gH�B�;~rxf*(�d��U�vԱD��{�.D�V0:n�CK�k83g��+�����+d+i��?�-���[�|���(
'���2Z��V�;�E^KcM��ҕ��|��i!�2��8x��H޶�i|��G
b����~:�1�of9�EV#�˟�?���.���o�1s���T�����}^8 {:�;�smFb��J�@
q�U�V����XVf�(�v�E,�Q1���N��(����v�E�p(F��eO��5e��˶c2\��/�~OzPEÇ��m�a<T�$Y�7`R��zX�q��&�c�vɨ�N��9o�[�ьG���Ӟ�>��#��4+8�yՌ�J�^�WV�[�cdf�������I��I�i�F:�A%���V�k��Ɩl�1R�#1�� U��ܻ��+is"�"�f"m��TQ�x����'�r�>O$�i����(wt�щF�˩�������%�%��
V��\O��r�Ʊ�po��Cv�:4�;�;r\ݩ����J2�	��0�h��
 ��{�%���O������Z�kV�É[��H|-_N���g��8�×gC(��/���=�G��L�\��w �n	 �H�$ą��f���b�Av�����ej(_�Qo<9�3�b�f�'��Y�2�%Wl�����ع<9D�VEJ�I��}��t[��dJfBxBky�����%��И{|y��#
� ����G�o9��h�m�@��9�#-}ϓD�w��+S�Z;�"�$w�G
Y�J��ʏV�+���lt漋,5�t`)P|,$6����P�cg�n��V����I�-@�U��]�{�Ë�2��F�B1���K�	D��w���o�u�vm��"�e<0��\�i-3	]� V��P|�p�$I=��
�N��;��L΍�8��:��o�1_�*C$��PF��Π�&)��u��s�=�M��W���=X>�䅲���v�LX��5���;��ǁᰰ�ºQ�4[T�)���@I[%����@���Ѫ�N���-�&8?(_�W��y����Z51���fH���$D��ƶֵ�F_a�<w�C��a�)<�pC����3>��=; LO�j�Ž��h��S���z��³�_���#u��x�e�b�䇎��R�9R+���5����H��w�:��l�����g��͋�2�7�sӰ��U�=+��� ��>3��S�BP�@��n��ͻ�xu�D�h80(�q���j����WBԊs��`�OQ�)��,�ّ��ke������}�\>��E��M{� pz��¾��}i�4�j�"O��O�bPf���d�-5p!<�R����H��1"�Q-�T�:�[t^�b�)!4j�C�����;����Or������M��Txӥ��k�@𒎰{����D�Ł�����' ن�8o6�>���:��%��W)y>�5�Q�B��w����DÒI1)�Fy�)G�r$*��r9M���^����q�|ps��d����������p��M�=j"����]!_E�F^y���y�݃�j�h��~Ûr[uaVb�����:ys59y"�d�zs^�"�1M�sxT?��%�Uzj
:{�ke�~:�؛�e���# ,} �2u�o}"�\Ɓ�ޜ{x�P �9�a��\���T���ߧ���z��xm�]��9��[l�Hԋ��� ��}��i,Z��f(�JH� ~�	nN���x�z�"�f1jF�s�K�\�y�uQ��\������o�/�Dd�I�4�+�� ��]�ב4�!W��"�`���v.��tq1�zy������I�N�}1������t�%}�/�,��Jqs[�a��B0$7���=6���fhŦ���ٻ��p��P�MZ<VpA�N�'xr�p8'\��5��V,׊����P����\�ST�.���+";�y�,�%;��%��w��%�c,���)o^�/~��Ҩ��O<�ZvGT��_��C{��v$����R�_�7���[*�S��f�Hl�0_�9|�@��jE)�c$���e��i������V���Y�uk�0"�'�V(���a�T{WB1�#ue�͖E౤W*+�\�p�G^5�J�3+}� ����CV�'�
�G}:�ds�m�#�l�{{f��j<���4Y�H+jo��ZY��,n��K����%Y���'l8��Ϧ���qN�lL�^�&��^*�;<�%�q�����Lփ��u�^��htKdQ���v�E��"�E��$�ݏ�*A���U�6S3oy�-r=k�Y�!�E��Y�	�^Q0����u��,_X�i9��yX�ьG����{��u�'Q������E�7�/&�9�:Q1��{�؜�W�$�w%���VI�Ed��p�����g�Ox[B������%��:�s�@�絞��Q����c�Ļp6*����1���U �-0��C��S�Hr���+g\�^��f^Q�?19�>�@;�0x!�}1�8Ѵ�x��#9�Hq�>�o�cD�Qȃ���+��J�l\vx�2��os�S.V|Jz/��8��5��1vU��S��-��~xq�X��+]��u,$�M��l�q��2f�3�&^4L��bpl
u6��XgJZ%��.��|~�q�2J����6%&��¨^�A�}S�Л`�Y�r^N�[KyrB�/GN�hhpH�e�W���+��_�%��ǘ#W�O}j}a��������y���Ulc��'�8|��'M��}���f��n'�x�P/�Ǡv7�Ytz��w�JD_�c�՗�{ƌ�w��u{�?�,nF���
$�W�s	c4�x��5!�%V�8f������ ��~g� l*����~� +��4�{��g3�7��X�C8��Y��.).���7	��A�U�zp�"&	��fƽj�9���z��ϡ��t�qNٟ�&U�j�����V��̑����,�P%�ڑ��D�\�e��C����9�U{��Fg��������(�k�t	 ���Qz2\^tmσ8#�dU�ի�FHBZ�X�eq�prv�=9SJg$$�.��r�,lV]�6�%ސy�����@¾���`�J01�7�I� 9����z�6��~2��$,�-]�O�����eW������tn�� #ܫďO֝r������Xnqv��(�j�����BMi��	�1���aZg^��6��E�Y&w}
�T�� 
&{;��������򈏴���Fm�!�S�A������(��Wz��ߘ�l��X�6Y���r��~��3�U_�C�:���47
�6�F�	�ʀ�����ϞI�巩l�oA���S��y��H�\n�R$�l���y���|��⣟��%e�]zx\�ؽq>�eC��[gF�ə�X�ڥ+�MP��|���"�Zd������|�������;��}��%�ʂwAEN�Je�g���m4[#���c�6ޝ�޻3��YڑdX�=����~�{>Ό�'�)���7��;�X���7,�hE⩐�c�e�o�aڟ<GK�E��0�ݟ
m{=�x�p�xt����&#X�h�����k��\]�ܹ�v\-�I��(�ڼ|6R\ &"v����W�C-�@�9�-O�#H�'@�`XOW�Du�$�< ���[=:�D�g|�=�lљ�[Tܼc��"D����:,�R8����n3���p���V�8�4�r����8��$E&)�4L����-o�^[Ae�n�
UtՃw7L[����$m"����wL���~�Pf�~�ʚ�Hկ��U��O������m���͔?m�֪���{������ͽQ��DUqeۑ���`lV�&n���`M*� ����IL$ĄB� ]�fh�N�2rd_�"���\���� �}��R�1r���V����W�����h��6L����w	������	��0�J��M��H�v
�_H"��cӀ<z�-ߖ3ţ�'@f�/E��ё����c��oz�7D�C�]����I�; �g�kF�[�-�����-��_��E�a򉺧+Mz����2Dnnݗ�~u��o3΋a.C�{�<�c�ݍ�:%�V��X��~1���2��X��Js5#S��RR�78�@( eX�9��>����0t�;�R��f����#������F�����?=�2E�.��+���H�}{wL����� �.{	y+TCw���������ʸ�.��^����֜Z�Ih��s�35IԎB�f�cm�67�6��!1�=�5��rN?�)���;�b���Ϯ���yn���!�j��>Ø�7���Y���T`��+/�A\�������5>��.B�@�Eo�EPm j��H{��6�iR���+H�+�nf,����M���!v|y[�pzNX���.h�[�h?�w9sB5&�#]��d��I 9�����3�q?�kH�*������[P�(�$�v�fo�b@ӭ���q�����0cl��i݊lG	/ף��#��3|�l����;�6��H	ʈ	�/��p�8����<W����FzunE�+%�!m^��4΃)B����y~�q��{V� �wdr>��J���2��̺X�?�a,ˉ��E@a�zt�SQ�^(�".����H"�}��A��+=�qu`K{޼���-��`�-�ƹ+�=K�PH�3��t��Xb�z�C�/W_h>Ж�ӵ����4��F$bq�#%�a׋�ғu;�N��J��r��?؛�Ŷ���!�?��M�C���A�Ii��J������>Ⱥ��3JH��W�y��9�}nx�k�} �2�F����4��BdT����cd�� �R67tRk!��>`Y`�;΁~���:"�oL�7�h�
y8" �~	];�M�,�^���^�a;��(Ć/�����hB�o�l��&����9�e09��ӮR�?��S���|���Xs�x5�:Bb��6�EF �L�DugW���7����SNCSۄ��u�ߟ�!���ْvu���U�\�B��zf��֕�Chᖩ�ގ�;�R%.0�]/�N�~G#��r
���l'��-�l�,[?�	(hDV1���� ���M<I3�۟]�
Ȯ���>�s�h2��FձC[oLB��'���iJ���o��� ��ً��:z1
�e���^{�I�{�X�
UU��o"䮊em#Og�O��[Z1�)U��7�V$��-�0}ҝ�mZ�����y)�K`�!�Y�b�-���a����5�zp�n�4Y3�T���!��V5I�kO��m�����qt?�ނ�N�孳�h�U ��Cl6�ؼ��Y�p�mW��FKR��)�_V�f"��1>Q/)ClD	�BuO`
�6C��P^��B����=��8��4�0b��7gc3���@u���҅ ���~5�����q�� Wm���e�b� i_��Wt����B��'��fĲ���XU�BXp�ץV�m}�̦�}�AX+:M>��X�̴?W/��}�$����Ӽ�y��W�F4=�'WH�h^�S]��x��C�X^-��r3�Q���^���o�x8�h��"b�  iN R��y�����MR�* R(W��G����I�Lv�t��=ʭ�m�ԵsÜ��5L60�^Z���
[�g��l	 ����_X�1D�����?��
�T���ʙ4_v3�c�f3��)?���ML�E�B���o���:���=\$��T�&����pѨ�d�?V�=o���|4X��H� �np��ka<����+���b*pp��w��Q��:�y��A�R�u=潪=̶�y0?�Σ�^ȘW<�R��=� �ݤ�"jY*��3Y�bF��Qmu�npɧHj�0��kA���S��U�|�<�E�о�6�<��6	7�h�˖�b��G]:�Xd�ص�$U���̫gJ�E?�k��5C�nDڡ�r��o*�g>�s��̯�J%]�����CN޴LW����BOP��b�� �{|��d�Lڣt�3���C���VO�\�"v���h\��ugd���:�����oE�%q8iL�x�a[�>G��=hXW���4�8�O�-���$f�u��X�ï�ϴ�a�UB���+撴�>ʺ�.��	�W
���k5�&����5e�U5���	���5�������'�<�%��@�\\����5l�=у�{���0�>�Y�
I��U�65�����w�%;Ւ��Y�z�v�SG���,1pK�v4�p�V����j��k�*5��KU�{tў��u���S<���a[�Guؿ�	~o^b�� ��W��A�F�f�>�;�_~OmA��P���ֽm�(|T�C+���7&�̣0�ޅ4D	>� d>S3N�m�h�+�;��͂U�fQ�u)���6!t
}��uf*	�� �SMh�>�1r�N��Qk�K�\�c�i�G	��ݩ��'�
*l$Joh����N~�¶j��Ã�2���g
,ܽ�]q��8y�������h��v���$��y�I�cd����;!az^
�7vb�z�ii����;��M.Y.j���bп����ҍ�-\���zg�\Q��#���3�iU��}���րT��ZyFƱ�ҹ� �ܚ#��B����%C	�{W{��4ݛ�^�V��?��j����F�S
;͘�Z�/�#��+_z�-��q��(�S	__P!%����&�N׎T{0 �ܟ��p��Td����0b�a�}�z���	�yZ������k����*�/ޥ`yd\WfW��6���lU0;d.��$_�:E��Y�]��P9�E��V��b��z�A�gi�zD-��~�P��	Cx�l��T���ϡ�=���{Q�'�[���i�3� ������ '6z�& �fj��/����Y;���hB{r�W���ۭ�EyBp~�ZИ�ߧ)G�~�䆂�j�`/�z��)�����h"�s��1��|~�~@�c<���s�[Lٔ}��߬�vx�p��S+Ŧ����7
�l%p�[��2?%�H��w��[(Qg|�ډ��7�|]�{�B�S�ax���1Vt�K�� J����üJ���Wn� ̆{��~>o�
����k.�0Њ<}~�j2�$'�qP�����X�M�]��_$�p��+F��\eQ�2@� ��#��u�m�%����Ŷ��]Y��Yx��]C�q�PGx�x@l��U�q_�d���e!\�Q��r�a���P����*���*�����k���~���-��I(ўLU�`˲�}k��.�I"��l~�mkSJ�,ʣ�#b >�1��!\�w���'DG�ɨe���ڧT�����{�V�Y�nvJ	3ة/[JTR���9�1�k����}(�Tf��BmY�Im G;����J�~ ��@ϢSx_l�y�~��{;Q�3@�@�GQi��6*q�������o<*8��� !2vW��US�����YU��u��g~�M��f	��*C.���Iˏ�ӫ0S����,<��܅QCGm(s6Q&O���7P��-y����� ݹ/��)mu8kD�y�<�-�s�U5�*���P�>������S��ԟd����M�<��v9�g�C'�QC5H����2=X��r�nȑ&�� �k,�X(YڔQ��$�PQ��¢G#�0��\2c�`q�p% ]�3q�k���[��&�<�R���5��&-��d$㈹����`y3k��߂��H��:�n����Y���1t)FD�y̔�Бը�����N������HSe��4�X��֣%�>^#��m�@Jh��70�/\v�ݶ�|���~r0��u[��Z�V� �DO����\HP�it�q%���@�K��f��4= ,�/����G����O�N�r��J����=៴��_c���'�[�z~.̭�MgLM�Qle+$=�n&#�A���^��Q���Y5c�( �ҽ��3���������XKI̾Ң|�#�j��Ta1�1"#���#{����P���,�s�s��V� :�����#a��y��^�8�������B�X�T��� +�EU�]x<�p�K�[Ou���0�����'!&3R�����!w����9�&���e���.��{�O;ʌ��R1Ab'Cu��;.��������BiC�o�|Z���^�:P���Jj�cqXd?���I�o:]��V�
3 �Or��	��T��[6�����҇�Y֜	->tIx�N����8����Y_��M#x���]�X��lT���7,3P���o~U�N��C�0��L��d����ᓧ7�)� ;1����7D-�p�+��{?MA��YoD.��5"�MqJ��xF���f��ŁJ��.S�{��I�O��`4�h��.�j�ޛJjΌ����d2��l�~�հ� ��˴�Bl����3��kj�&L��;qd�c���x?kt��̹0��I�����e���N�����s�л�N�(��ٳ\��),5V��������ʆO��6��yl�[]^�|�ӔK�V3��ӣ	���͠�ì��k�Q���AI�6�(h	��<ᘍ��q�g�l�7�N7�M����%%�7�3E
�� ~�+�hH������:l��A�k�!/������#A�ж\)��A͟b4@��U%jS���#a�a+T�3�F�ځaM��ew-̲�K����3{��k�wb��2*:��8ߕ���D]c8|�u"����
ܡ����� �N�qC�� r�����Φ�V�[$T���� ��㘧����h/�98;sw4�hY�Y�ߔ�_���=	-)RR[˅f���Ok�
�xt2v�ߵw-��_��z���虲Z�"��*D�ih�ϡHt�YW�=w�Z�d1[�,e����A�#����V����&ŏʋ��"$���/�>��
�Q�� �[k	��
J�{�q�뤣K��'���jh�"�3�q�jÈ	��+X��W�'���QB�R��c���4ǝ�;� -`���|32��	Wi�>#��.�$�]�/	�b��/@֮+�WX�l4���t>�hQ�����ox�~��1
W�D�a�}�����>#�5�z�*Ä�Y�@<+_4$��i�)�(��*DУ�j�ofofz��v��F/��=1}�s�xL�t�t���P�M��qM��>t���e�	�����R�ky�Ŵ�uZ;V����	��m�H�^�.fJ���I��a>���?\G���M��2���U�x���/ԐE���ߠ��m`�r4�2�?0��t�����zU?�LOB�32���r���T�ъ~��s����b��K�4�H��Js[,-��iϚ���df�ՒU�G�|��c���b��6��KK�N������3n��PlK�3�:�,�H��W��'eEP�#cYS�3}Cd�Y��kM��4�!���a!��d��U��=J_ذn�M��D�ON���!�lo�,;��ΛE�����/��f��P�-,����=�iHw���{ɼ>�H�:~�����=i���Z`���X}�A?�]�	��y��`�Iڟ����P��DJ~��7��5���%D��V<�c�5�J����d��O$_�xd4XYj&�}�����䍜����u&&@�S����U�M5N��*w^�̶}����A�`��ps����݉��o9�uU1�l��7f�d���a$��X�ڏ+���:q4y�D�I���/A��x%T*�^�~�&�P`7�������(?��oX��j����
��4�۸�y=�zƾ��d�X�Mj��)-������Kgd)���o$If���^s��vb�dk���+E��7�'z�	�� �,4IzWz���NW�w�I0sSБ^km`������x�ˤЄ�y��&��6��*�\ �3t��f�m�K,��_�	S*�V~b�T�z}�Q���r�[a���N��R�������G�O�%B�o���ffܲ����ÉȆ0h+MW'o7�N��է��]}��hjύ$|��^XX ��5��0B�us�ky��O� �P��>����Y)T�O�[����]���d����;x>�Y�/�fک=
