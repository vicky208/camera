��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�U�X׶�C�w�	��������m�	T��a�m�4��:PR��/e{ؼ�6.��\��re79�oѡ�40����pg��`��a3�`MG^�5���bc5,\n�aT���F"o�
rO����x��ٛR��֎��0���)�Т���q����Bf ��G��Y�8.!觔+�m`��0�+�T0|ώ��I.}��bUp/��Y-0���$��kI��ᖢc���5a�e����hN'����C��gkWaXeԬ��= 2t��Bx�������:DzX�bF/�H����w����A������(�W�4�W�(��j
��@#��7z�ñ�+�ҿ�+@i��ֈ ��z����Qt�~������`���2�S�^ Ь3��,��x܎(��umZ�"¡E��,�
�$�񅁽�|i�10ˑ=�S��b#�H�F���9�~����q����]s?��%��(\���SȇdmCV0}A��s�]�sn�c��~Q�m�#��e��jdB��;!��31��F�7%�����m���*����X���"D�q��!qۗ|H��7���Bđ@Y�qH�R�H�����B���$,P�F��[LoƱ2d�Ϯ�;�MU8�S�D�̺Lq�kӓ��l\�ȣ	\>y��g�G��|�\��� �[�RT\ށ3kf�N��>
V��Q�*W�e��֥� ��Ky�������h�hE"L���ob��R�d�w\g����)�yk��(	��epĈ ��]�{5(�����H,慜_�:P+=�C/��m>�%�{-��H�"}>��J��Z���Y?Vb�s�U$`�w�U<p�n��"�Q'�!��@����z3��ץ�k�\L ���~�9	�H���W�R۴��z�h�H��]�\�#�d���t'�����OTJY����i �m���4NS�?�s��3�u̦���nk�$�of*���D�X ��){x`
�O�x?3�� ���[
=��z0��X�[�����,��_��W|æ�G�=��"g�֧�}�6H]Q�>�T;�R��"�� U,p2�fFb-�ϐ��#S�&���`����\�e�v�_����ٱ)e���U9�*��ߛ��	X��ӄx70�z�N�So�@���~Pݺ�>���?sF�~4��hSP?�9'��>F;�nM�eZ	�����t��9ÏT��"ϧ��\)t�&L�[�}���<�����c����h���Rs��fykB�C�|���{��rזV1蕆��?�2��l�k 8����i�` 	ɞ!Y�$�
���g/W�8�����C4��I�``�mC����'�cA�/�Zӌ�Gm�'f�p�s9m���������_�dz��2�"�'����`�ob�lF�jo�v\Au��y⛖���!g�E_����	��I5�.r�����x?���ԣ�P�İ����߄��yQ���>1�C/N@�C��,q�7�?��7�B�x�Տ���M�7�����?:�C�Gߟ1�ɪ��%���Dy+ࣽwJ؟Ɏ6sZ-�������6��q	(�����ˀ7�,(:�a�n�(M���y��hx�����w�x&־�����aǳ��	p�%Ő�g+<:)	����Zs�OL�(�e�=F��k��'�!ʪ10�ztE��t��o��`c��������H�-1����(���(�^�x�K�v�H!Ly��o-@3���h�� �V?L)�a�k�q���z�T�:-��Zf(WB6�6�(`��4KA��i]@��M���U�"ũ��|cд NTc�!h̀��V��^�aV7Ÿ7܁w������(��١���励4�a�l<F3t�O`)��.��Ae��]ɪ'���I�#�����u؈��\M����g�ٛ��ҝ�#e��Kk"�����=Ĵզ�2�*���B[0�Tˁ_�INC���(��'�
����Gl� m�D�Y�EP�w�"�p�k3��������u�A!��6��������|%�qJ	M��� K���`�go)�Gdq���U�]xçeb]K	���b�ɧZh���;�����Ǥ���C���R�U^� r���kg�*�.$<���|z.5Юm���ȓ7�΃�f�-�#�jԲB�{!�)��`p�!h�t�Y��S�N�,6t.�����d-���ؼR�у��6�L%���Bk��g\#Q�5�aaBH�Uo���:e�U�O���]��#>�ӗ<�i%~��t1��E$VK�)]T�F�>0�r����W"�6VY2$UT��K��!a9#O�9��[�9�~���-r���j���7�V��h�]���g�9��|W��&��%$<�\6�V��ޣ�~VC��5{���Ш����{EA��zA� ;�H���C)�
ͯ��V�₰*&"�+����D�W��Cf�2ݦ�}˺,�j���Jsn���K^$p2���id�^cj",� B��S$���=�i��K����\�CY=����*�0)�d����S�S�Z2�m��ɽ���g��$&tx��(6): jRu܌oK_���6P�	�F���s7izUe1:DOiȶ����4Ii���>�Ie��}���.I�.g[�z�y��j���Q�xk���=��=����i|m�A`�R%���k�R@	�g�@�)�ӵl8P�O����Hc�ia4����A�{gol�]b-� e!O��򹙽�)�)sP+|X칚	�]��)-YW�g]�KA<"�:�������AO4�m�*��9��V�t�1!ZӘ9�,�<�ƈy�|(�t?
���H��k� �/���D0���AZ?i~п�So����+�\v�u^f�G��5�c�rJ�H�R�3��R�z�Tl�\����|�zЄ����9�Đ&��শ���k����=f���1��#g�Tw\9�"�rG'm�	ԹR�鄮�D���i!��C��p3k���j<tO��H��/�ˊ�At���+��y�h�H$X�/6S~P����
�67��	��$�&���!��u�m#�XU��bʦ[�AtU�+f�Ε�(|åR�N�qՠJYXnocc	`�����ɒ����l����Ϧ�c@����3����f:��a�I3�7�����w������£�)f|��,Z�7�w	m��![���x�<i3�I^�v�Uɑ�u�LV7�;rp���!D���zj���hD�[��H�%���ǰ̰QÉʟ�>*yG��U�SL��oM�xB����w��7�E��<��N�uťwЂ���*�LC��: ���q���28�/���/��_R�aE�뚢�A�ַ���N,~��ҭ~T�֬ͤ.�L����h�/Yo�_�ݏo�%�e;>M��*g"ȗ��UwSulz�����?6t@�����J����C����+p6rl/ZSb?�j�w{�I5PkO^�A�u���ө1��d���'���[�6:?��G/f!��R�� h)zi	�"K�A���$���g���(�O�u�S1�@6�/4�S��� ���!�ƶTSq�t�����;�7�)-0!�X��ܢ���P����d���_��K//T5a�/+��\!%CI�x�y&<<BO�P�+x��(6��W!�.���%���,�w�Tz}��z���]�'���o1�X�W9H%�vTP��v
R7���&�h��
G���»�7� �y.�2_��
 ���~Z�3z���Z���32ZzN9�F��F ���>��x��$��w ��+X����n�YG����K�7q��L��ܪ�:8����"���2�U�W�_�K;�����b���a�d�3�/�$S���u���.��Pry���д���.1[2���Ҧ)b;qk��,��/1��3�H��-�a�zȕ]�ođ5�6�/�o'���z�l��o?0��J�	i}�Tք�+�_R��d�{�ǡ_q��&���,񤯽Le��w�F���c��.X������� ������}	G��k�N���7R��e]��`#��3�+��l��(�ŷ�r[�� B�IUƙ�4E�j�_D8Y�^���>����B��B���΅�iR>����Ax2����qf��4VT�r�*��-���m�]a�H\�<�CS�j�\V<h����ÄTM,ܷ�0F:(�����O�I�\3i�Nyr~�9��s؏8�nrԣ����NjI�v���:�ÓO�F�����V�V���d%&w{��X�I��)]1�1<��p�5f��Qk�e����W�����V�K�>(���~I��Cb{�y�N��_�pg��&�����Q�]1	Ѵ�}_������Lд�z� �v*����3N�e;�۔w��H�f%�z���I��PS}iH;ذ�7�k�Em��W�}�N=���i���X_�1��&��&tl�Br�i��sZ��ji�=4�GP�4���nM�̍ q覆��>�zTX�����t��cXW�D��[Mٍ�J�VS=�dJE�Mf5;P <�'����k���{���H-��4���<��ݻp���H1�f�g�(>Kml
2tS~GS�[�fAkf��"�ɥ�"����(L�ǟߛ-����^! OK�����h^kۑ!���T�)q�0�Os��͏�$����x� �*�|:�̹Ç8�,����O}y���dop�����/��'5Eо�p�E�M%��Do��\�w�m@�^
�!�����a}�$�G'
$yտ��}�LvN�->��X"oSѦ �=�cx��|��U�d�p|O�'hi�B��3�Sc����2K�k�i�@ί4/�y��=�w�8����WJ��9S�晱�D4�L��x��{y�NŇ�R��D���>Z�_���PH�щ`?�N�S��P������_ݑ���[��HP�-���C���)�>�
Y^�X�-�Gz<Zz1"�H�!IX/B��)�������ˉ�����ˑ�:7�p�X+煟��z�����Kɗ|A��<}3y�."կ�>9�"L�I��A{�@�Nn���,�(�ӱcH�*��	S+	\FI�)�'<���"+���w�9f��5#�0�f@c����b�"G��Ǉ��5�NмU�*����c�"U�x���%6��`�p�Xqd�K�|Ye�"t���iȘ���u�g�<�2�����'�Z����Pb��?Sy�~��^����I���O��b�
n�/")?wƃӮfïL��_�d��d:l�F1�Uӻ D�>~T=7�N�g��VnX�GW� ��ޢ��;<rn�Y4��2*Mƀ�O���n�� �������g��:FjM�t����G8_�;.�3�B&e/u�y���I�6��w��g�o�>�-Z�U�w��G�Q}{��If@���r`�����d+UUY+�%�g�ە�B=\X�bణ�����,X6��L���ך�)[�Cq�dL(�0��9�h�DRk�bߙ֒����bwE=����wNM���)P�2���r�����|z�
��/��f�l��iyB�8C՜%~�bS��
�B�2d���}.�Χ���P��o�e����{��a�)|�tb�҆�$VQ��g#"��7!�e�e�Wf�[�[�e����%Mu�����}a-�YdYr�&d�l5�%,��o��̸�C���X7pトa߻�k�n�.�ow���G�!�$�C]/E^�ff4:���E��R��\.�W 9��8㜝܋�{5�|Ɛ-���+�"�E��+�Y��	2��9Z����^K.xq��s?K$tF*��W��BI� q[iA�
w�{�nʝ�!�Q�d5���9�(sg
/���ks���ԫxV �y8�Ct2���O�b�_VE�^��<x��<����S��V��D�_�l)��Ɂ�����̎hê��	vR�Ĳ�	�%�m�:x� {�K��b���ns<+�U�
�nٸ�n('�1Í���󻡏�Ř������.��kB�}����#ݷtu��2�Pu_;"!���=�w~I�{���prN����D����"TY-��Z�,M�{�^D���p-����k�^�Q����|��~Y1�=}�*4t����K��-Ж����LT�H�vė����9��-����̢�嵵<�Dݺ}��҉u��$p��^az��k��ᨺZ��J�{��]��j��X��xĲ:�%�l���mB}��s�Tݨ�\XX��_�'��	Еy����Ã��ˊ}��I
f��W�E���韦���'�[��<V�m�wI������K���P�	��,1�.�f�9���58��x�|'WƤS�Z�1ڴ(b[���^�+��86����ܬ&4dV�䪀舵������o"����q8��`ԖN-��d!)d=Vz���> :�K�c��1���Ν6Z�Y?��X���$�G>���!{
��P���uj_L�:	���[�}i��o�;%9\p
"Udf�I?�P۶\�o�tR��/��&u$��FQ�PL��R?�[H��j�zrO�V�c�S�	�����}0'p=��gYu�.�;Z�����~�TO��<?�(|[aʔ��4��#��E�,��r��h�ۃ��K�ǈb�?yX2��bD���qczX�7@<M��Y{��ή������L���j��Y�'�LrA��.���3�c�as��8�n��ye]n���=$dŵ�����Tx:+�*n�l����ʥW~��e����\�鸆��4�Z��D~�`�٧�1�g\k�V�$�a?܆%K�����yM�	�#Lb}i�d��B��½j�<��j���ae�q�gΰ�L��?q;
v�k'���K���R��jVzNq,�-�:�7��G���/���۞�.3�_�Y�0�-ݹ��R���'rh�����gY1���Zg�	��,�V�P��ݠ�X�4��h ����FkO&�c���G�C��M�j�IQUx�mWJ�x��Vd���[wC�������i����'�<�i��LzAOd�">��n.d�NSn�������NDfC���ze?�C������.'L��>\�ϺQ��qZ$}�!t;#��wV0�*�a�FC������C&����$��k���L�7y��<:��=��OU� 9�2e�J����{3T̪M�IVD�JY�Fs`�Ɩ��C�n�ki�D6�=�'�È�.,;��}�����^�݀8�O�]����JO��Ԝ{���/v�a��a�R��߱��!��J �B}O�7�=��ѳ�1ߝ�m*��B�xlw��S�LQ�T�3���_$&��)����R~�n]ER���