��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V�B��&�8D�o��t�� '3��r+-@��
vE���Q�Yn��+���,��f�h�]�Ĥ�_X*E��̞?�<tO� y�3J8w�_/x\�2Q-W�X\S��Z���kr�N�}iQs��a�����U���<U�;+��a����s�[Ȗ^Z���Sg9�쳉���'G����$��<�]\�ۏ�xt��M����g-`�-S/���[��H�:V��˄\�C����PuMu���''�ڗ�)f�说��/2�Pr['���g+f7�F�խ��k�]��xdD}����7
�W�D��P�,���f��?΅4��&�cա&ʻ&�6�#i8�Ϡ_��r"����V�c��߽�d��U�i33��Mr�ܑs�̲�Mdd�cNա�˝�0>�4��;E��+���[��DŤ�Bx%�F#��ĵ\�M�j��z��}+�1�͊=(�'�e�EL���N��Ae�ܧ�h];6?m�9��݉�(���%��NLo?Oՠn��t��0�v��`ga$�r�\Y�l�wI�u�	8��CMa����8I�Hh��w=����}���k^�!Ll��ha��؆zX"pE��i�\a�u���-��ㄅ�<UD��ҥ�@V)o�f�+���*����ϝ�)I��� ��/"<G��&��}~Z~{_����0��
�i��Y	.��X=��f�j��-vy"V�.=x�[��IƧȩ�����pv�4v�&��gq��VA�W�������[c�t�X"To�N��3�����ed��`�)��z��	 �hgN�A���5�si�
�~�f��c+��6��&�{�y^v���ev�J�}��r9eH=�E>�ˤa�64zU�b4�P����/�P�4PP����frIh2���1�K�pq�g��t6`|&���@fT7�	}�0���c�X^���wr�d*+�ϷamV��h�bI�1!��S9���~zF��xE)s,{c�5]��4rM�G�F-�=��x�@���_R�:����+y���B/@�(�Ck��
�������c�s�1���$��W�y�����4��������v5Ja�q��cP��:G�����*���/aMO���ʯF�ű��?E����;E�0e�Z���@�-"�yW^O(�����K0Ix]��~;��㼍��� =J2v�"�Q������_D�"7be���ǖ�Fz㎶֥؂��BĦ��O�-�P��qq�n�b1gB�.��ܣ ���jH���k�z^U�����]`�tu��k�&���~��ֈ.ښ�k��G��O������S���"ɦ��A�b
�:�=Tf+p ��3��)K:@�]z�x��=U慾�6d"&�-Qv����\|�^��J/�*�������)ĉ�{�����Άs���!+z��9g��9��vo7�����R��Jgj�@+v`Lb���r�/aS����̀�.R����b�CF̱]�'�M��@I P������s��:l��HX�n�QS�R1-Y$�^��� J�l�UC�	Ҩ����*xL�NdR�������C������3��f'X���냎�
������C�����D&b�3�0�}���L;�@z}h)�5��U�/�_�q*p.�ԕ9,U�t壚ht:�Yx���^�g��K"�9�`]�Z�hkt?SW�yj]�p��e|��+�#�pz��߱Pa`>��}���31�w��b��5��ǩ��Yy���Z+!R�gJ��.�m��C�]�Ij=�� L�3%�����G-ۨ.��:[�*�q�kf��0��K����y���a���wg�(��z$�5�\�Y$�7�T�1�=x&5�o�zZ���P���-!k�������, *u!��w3���,=1˾�h���tk�նsٱ�x�УJ�ӊ��%�Ф��"f+c�̙��9 F��n�zJT�Az�W=7&�f2G����;��b�	R+��1�G,�2�ٿ�b��Ej_@��d�#}�>����>�?7�=y6�cs�4�2�jaR���@�Ai���~��Գ��h�ui0FaSWƎ�L�� �&�8��X���������:9kK������'W9�|�ZkA���ؒ�1�
>q��`L�$�c�72ؒ��Ο�;�O��а����s���I��}/�;�1�����]���o���'ڕ�i�M;�{��Xrxz6�6�_����y�+��w�yp���J������)�;���\��`�/��T(�2>7����!��C�X�Sh�mLC\�Lf���:�y+��3�,ӄ�z��=�n�f�"�#&頎1^��H@���2#l���(�dz����	*�		��P��4ߺ���\���f�T�!Gqa���FT��h������R�������n`k]�]>=c�Oו˵��}����/N�	�����-E5xŇ���9e��Y![�����?���Y�n��x�'�X���'�߫9�t嘲����c�t݅�=�� ���Q1r��8����k�ߖN�1��!�^�7$ �z6x<�d=��{�p�-B������d�r���H~ ��%(���ZU�[o�c�Owt�"^E;�ii��l뜅V� <	5�����Iט�Y}5�W�HSO�@��r�;R���<�`T���҆�}J7����01�f]P�+�Ҿ)+�i�u�������5u����n��Y\͵��`b�/�$���/.n��/R �!(�ƺR#��	]�uGp�0�����O�枰/���, �y���ڠ��Y+pgS�� d	�0��p�ȿV���%��фh�`�0r9:Hn����K�Fo+䝕�>�������:{Q���M�W5v�s3��5�K���O7�N��W�`�ћu4?�����Z����)Zb [o���ok�x���N*�um-�8���
�iw�S��/���|�)!q� �:�閕�x��єq�X�	�X�60���/�VR��.2�Ϥ��xi"�i>oԽ��g��\Ճ�+8�oYՈM� U���>�C��x���܃5)��)���p�����W���8�3T���`*�z@�c7L9�c[����1xSf)��*~k�F��C��H"�L#����*' �/����s �}��`'���0���X�l4L_2<h��TZ/R1�����w��(C����b,�@\������z��v3�'ՑC�(�����d����v.^e뙓a^�Jј��i<o4�E#>���3:j�lY(j��VP^��e�1([�� ��(��}�`^FW�v�\��"�C���g���[g���GDI.ݶA��S�p�wq�f3��l�Q��-na<�v� h6�}��ՠ��P��W�j������υz���D��_�p��=�"���L�����Y���R��m ]O5�"�10�!�wA�� ��2��1Տ&(�6��*�-�}����c���Za�R�(�{nx�]�=���7������*c�Ϳ�z�Z�qC�}�s��哖��j�ig �v���3�M�q_�B��.�}t�.�X�( ��1��̧i�@�s~�u	C�j� ��!�y^��H�)�^La٭�e8��	Z�r>�`��,���U�ɅØ�V	�O�q�oYc�RԸx���� 
-v�diFxͦ���zr����͔<���:.�&�����7�g���'E����T���<�r|'���]�׼��W� ���k�!њI_�-���(���4�L?wP2�����-tS��z�O�D;j�+��P�TY�
����~!ycرDw,�ۻd����Z�7�Bt�ԛ���k"�҃T��tZZ�OD8C�� ��a1C.��7Z��m/�|C�!Ş�~���yÎ*!�u�r�W���7`�|��q�k��#h14�
��<���"S�$~��ɉ��Gn/�l��VSweva�W�3I���4Zw��؀�1�¿o�wB˅�F}��J�6l�%g�,�����E�o��n���7�	6�j��)�� xɕh�����m��j-Bm啯��$�����}��(Ce<��K������W(�ǳ:�$o�T�%%gzo�^�g7�Z��;���u�r �p�����f�b/J7�:0��6��J���y��o(�{|ː�I��O����|������(�|�&�����5`��c�,X/�/�+\o�z�s���k�cuOy��Ȝ��_M��@�H"d��m9?p��}�{+D��q1��7zΕ7��lO�T�� ©�|&��>��5(��+ݜH���0�G�g�^f 8��Y��%3vUѻ׫�t3z��߷.�r�ك�wo(?5_�4n�M���
��z'��d:|a�2�U>�~Ct��M?J4�$�2A�����n_ηw�,2��l'$�^ʌ��:���.i"���jN�O���"q� P�3S��(� ����TP3�;C����S}>6压����!��x��~1�H��W��p+}�|j�:G�[�7�Q�a:t��YT���R1���`��H�k�:�q�.��-�C���DĈd��M� �h�8��.�
b���^{�ub�vI���wk؜���'�-)i�:��g�|�bÅ�{�8d(U ���x/)���>�y
�Vz�ri�f��	=EwDR���"���zN�\o��}'�e���h`Ѫ)��-#�oA�'��w��� M���go�U�8�h�C�R0��t��=�et�C�poGk}*�h�i��Zpe<|]W��P�B�{�tD�x�%�r�Ө�Q�Pn�p�~\=�'��m�aD#�pT�g��s�e&��(�	D��K�����-dЗ��]Q�gx��n��u��y�iZѵ��º��n�`!����G�E�	�A�P���������6%`7�|����+'��.�h�z��B�x��DlI�-lXۺ���l$�mEh�0<���p3l��ڐ��F���'��yl���٪���Ž/֯� 
e���Z���$s�w�ۡ�jO���BG_���O3�=Z/=ҡ!DQ�n�o�s�O��"��gk,pEs��z���tt0��wۊ�&0r���
fN�X�漳,���,���%"Ħ��˃ \���?^���Ef1@�)��4�����R���}�W����=Y^�#�6C8X���Vu�3���m����[���A>O��jI�Ć̏P�^��:4/�i�s����6\�OCA+����XP�3��������<
<}kuMxP�k�ǆ"�k~���r����y���RՑ��ړO>uh7Q	��-I#jPn�HY~	��B���������<�N~H�b�4m���ق���Ň��.���zy�ñ4���X�k.  P�����Wt����&�o����+N�|۫�/�jR�'�H:�^.$-=��(�_�����'Y��J˂>���H;R��񦭐s�AV+-�)y�4��
g�7Qv�wN�������U%�q0���py�]sq`�`>yX7b�?��~�,K�<�.�Y�/:;���l�և�6'��+���L��:)��Q�J��d�TH�6j��P�:<��@5��;���1���ӗkT�Bw [����m���JO��+z�O@D�x��9�\�!ɒ�7�$��E���'z������	��&>(>�w>���A�*��+�X����)}9qw����\�֘�=����#�xHR+�T}"ӹcFj��k/`H�=�V�8�n��Ey��,�rn��5t��J
E�I1�8�L3������%�������	Zz �jU�qZ��F9�jlTwv[����@���x��N&k]���B���#�ܬS�|T�e��8�X�q�4rw�Xk���~��=���g#�ǚ�"]����������w�T�9�v�h��E�x�eP��z˥ A?Y��'�}C�T�
�q���sG�~�o ���8x�=e�bB1t�\�������tc)��;��h.V�ծ�9Ko6��=��q�` ]��AfdЍ�Y�l+�bUݾ�j����F<|��[p�-�JL�W],ŏ����H�`ʿI��ļ���q�x/<�L�}��c�)����j�刖NU����G����[W����`�yyͰxҌK�D&r����I5o�T(Q��x�c�)��3�0i=�n��R]�<���WT��l�qr���NiDX��͖w�C4���"?���<E�V3��%[y�M����^'ɏ��ò�F���>oNюf�vwp���$=Q|J�X�Di��D-��b����n�a�f'��Z�-���r����E�����obo�bnc~@X�GT���u��Km�_g���
=o��V#����;K�~�F`#�H�-��!��M2���`���~��V���Uy[�į��S	e�'Ed���jI����?�~Wg9H)�3�lXB�t?;\�+:A_��vW/i64�td���Elc�ل�>#�"��R��R�j,�_���#Ã=[;�o6۰^vS����:|<��l�E$UAV>R1!L�٨q�e��Rqꔺ���%7�vri�:�o%mWrI@���K�T?Oi�jV�2.F	��z�v���0)�������X�����S�u6��W��]�� �{=�IL@�O �B�[p9�6��o�2�w��	#����]��M���2*�3ux	U�9���Ҵl%�2���/!��(��§��"vΚ�ݓ�+�܃d�k��<�oCį�h1SR�Bk.N1��3���yQ��vִ�V��J����X��Iɴ3����c��f��$�%;�ݘ ����Y�~Ɔ~C7e-v��W�cC�81�7��L�o_�����d��߲a�Mbm%���$��nF*s�y��	.�Su��\�ݚ��rKl4A��q�5�pT�KL� U��V?F �%w��_*ì��������t�E��(�"g^�����tc�0�i2�>}�ȍ��N�b��W���-[xӀx�r҂���I��0EFdJ���-k{u�=k9#���M}�޹s7u��ɩ渣�Ɗz��h�XAe������8f���ҒM$`GT�������g��|�L��;���#q��3R�q�"����zD�?bx�e�P�l�3Ē��{V�3<k��
tT�9�H�.�[=��G�P���;#,�fq��esdӎ�7���O��u��%fʸ$��xX��M[�4�XCF�l˝��Ml�"U�;n�l�N�Ť��sa�~���x0��^a)(B�E�@���kFz�/��R��2Г�����3��0�ت�پ�$���7�˓��&]�hυ��Hn��YD��N��Rh&�D�%����L �fl ڋF�Ҕr��q�"�vj������qRI�Ԝ��æ"v��i���N�̦�f�s���˃�֌(���Ln*�5^F⢽Q��#n����iԕ�2a�%hAp�P���Z.�P�깫l��Y�:p�p2{m���0Շ�^��\�(�X���?f��NI�����:���đB��;���YI����`Vc���o�tbu����6��j@�I���:r�8�y`���oD��40Sk�Q�ȴ����|�5M�"h�.Q�S��p�����ۇ0��#���ti�8>8*����V�лO��hl�?�,�Y���k���Jz���R����g3GRw�n�ۂ��2�������5�>� Lw��1Z�aZ��a���6��v��Y��(�F X��I�f�x��>�'ʮx{B�c~[�*BX�r=ʦe`��~G�d���ڤR�t=�G��ӥc��
�ۭ���h�(8M�"8�ǂ�8ד���Ħ_k��e��KM�w�,i[��]�cc�Z�\y� l,�A}vLpL��
��H��UKڀ���VM�x�т$Kr�W�6�o�_[ʔ��w�<��D�,�q�]���� ���Xi���}s�=%&��r�����*���ȍ%P��2Ujt(3��T[�My��x[�Y��u.c����`~�qB_1�І��>Eo��èI/Rڅ�e����b�d��'g3�=4��b��'�^2В^'�W�>Dof�Ǚ�(���R�^��kF�s6P)�w��ۡt�9�sB�����Y�sj�)�ŷj�Ae���cT-��B�����D�q��� �gt0g���v�#Z� �xJ)���oP�q �7x��="t��d�Dޓ~��pE��X��f]��i-�+�"%S+�ϫ}z�\�q����D��M�1'�[y��F���Kr ��?uh?����!��������Tv���bVd4I-���Xs$�Rq�F5����Gn;G����Gp�2��Й���S����8��iS7���T��*�HNk���YC]8/���m��{�[@'[v��43�[��#nè��:1���\�S��7��i��oQ��	t�$���V�Wx=ȷJ���.�,�9�ބd6?�}9'WAჟz�|�|����Ȅ��e%AL�j7)E(H����աP�qx����q�}�Rb�Ω�u�"�T
S�)�/�"	x�y�,�U.i��A���m��B�u=d�s^�A��6��b=�dy���c�G4N�>�Z7�*B�Vl�$���N&���ȩh�b��_�����a� ��U�sp�W/�����\�Z�~������(�O��'p4D=7H/{���ϸU�U��|��u�WrB������M˿���AYeB|_�@	�Ÿ�$<�؎i���R�.~�T�<
��u�xf�-d�3R�����@�جŬ�S�c������xzi��魁�Fc��eѢ�v�����3P����`��ui�}Q�����k�"q�$�$��ᬭ��3E�*![�g��'-��N��gFқ����?���d��c��8�(�U!�PD;ea��! ����	A�3[2�-�������ܿ��"���~��皅n��%��~�#��4�7��l#&�����[�����
�_ij����CU�����Z�Am��x1�MX�:��u�;{χ�����w��[=�]�8�մ�u��;�p�y!��g?+��E�Εy�s���u9�x�.���ts͐�� ��0d*Ë��|��`�15�0q�bN�ɷ�k������W�"O�f��\�{���������i����e:�5f�׾��A0���F,E�w�
$�0OKP�l�Î���f�Ї%R���Gu�s:�"��o��7T��ijf���>�n���L <j�@SIE�zWdW���� �	��^Z��t^���`�"Ӻڈ���w�5p�f�hw���j�;���3�����1�%4,F�m.����,k۾Ųƹ�υ�3���Qj�O:x�Qϝ<
�E�=u��C��\��S���i�� �C�@;�k�`��y�͘
KI{����{(3�r��G;f3�䳌��8Xv�.��d|��gƥҭ)�tA$W[yfy�N�	 ���1l�L{�W�ɫ�&D_���f�1jڇ9�crg�˓�#��<��^ �X"@�
�_�ꪙ��`�)�GDY �odt^�y�7�X}��~�J�$����l,������]�d1 ^lO�;p��%�8t������'�<�n*{4����z����Kڧ��raL4�4;㾊��~�x;�����v��F��_�p�U sD��Ks�S�.�*�,�3�q�x��V��g�׽2��$�o ʺZ�^1�NՊ���D{"��z���|h�u�R��*v�� �&z�rIu tR�}�c���� a�d�I#�̝�a�������?	O{�F�j�&/��?83�k���7{t,)���R��� B����v+y�ނ�K��劍��q!�\足� 7%	�̼І|�'���Ulwra!�P��/m�ӗ���T�M?����a��0k��AuOZO�i�lgί&�����O�fl�#��/?����׊�~�~��/�ŕ�^��r�8��׌�:(�ۗo�#�e�������]�_�];��'�y��@��5pl���y�r_kف�XA�[f[���h��4��t{����߇��E�Y<�Y�g�gi�]Zh��Z�Ú�o��l�5�[FV��@s8��'�	ש���@c��4b�=��������}Á�6�oC���
G������g�'�1 .<zG�|S���ܖ�|9�inY9��i)0��!��C�D(�&��e�(�5�ˎ�}��ǩ�H�G�����;�^ai��č��: ��� �ǚJ�T}�gk�i�x)����|�?1>챋���)H�3�V�$~�܉�a��;G�ۖ}����;�R*!O��}D	\��#D�c{�/�d�B���D6x������y�HD������Z�:���1����!��Q�)��Ms�Md
\<O<�D0���q]7�f�k�5b~,�E����iV�2�����=D*��k*2� B ��z���0_�������'��W�02�Jv��n3�K'��~�a��L�ǘ]�YW��?���']�[)��ܬM�3R�����שb.]m��˾HZ���m��T ��zs�@�R��Ҥstr�pe�t:��5�C,�68-���Ao��$�7kh����?��G�@�>|��N�Qk�FR��u���Sd��+:�S�/�X�jvMX�T2ϊ�v3p���r�eW!x�Z�9� b'�~]��c0_J0��x"	&D�"���� �LB�Fq�T'i۵
Ҥ��]�����=� 1]o�V�W�����J$j�J��W�� ��(eĽ=s�A,�i�B�-u�	��n�:M'`J��n���ʘ@d�{(��;3	��g!��# �\���؅��f��������/�!W�1d? �Q�x8���m_d����/��Bś���(YjU�x�o�=)1` CP�2�a��b���z(VΤD�G�|-wٶ�;_c��
�pTNrC�0L=<Y����#4�/k�q�= 7O�/��{u�Ľ����W��y �\�N�F̠?���TUb���9v�e���=��Q)�������ޝ\y�Ӄ,��`yʇAA;�K
U=�z�&X�9v��J�{�_�
ٓ��EL_D�?{Y�<��#Y��D(&!�K?��nS@p�Qog8(�3*��1�v�:@�k�� kd{�hnd��g~���y��	��|��F͌ ��<��M��vr{x��8w�V�̗γ�뉈^W<�a��(�$Q9���Z�����ew�}~�̔(b�ęS!d[�1��`��/&���f��R�P�pss��5�d�8�'��2�yx�A�d��k�&�a�SߡP,t�Y�h�����z>R��T^��#��p��iG�L��Nv������dzqB�P��-3�c� �r����W3h3���/�M^��&\�-M7D9��[h��P83����ʵ |K�o��)�L�#N�������Ӈ�W�i�OME���ݫ2���P�uWj^�h-��p�3���p��Ou9HP����G�7�6>��/���I���L4�-�1*�l&e�ㆡ~����v�dU{ �dAĤN���)哗���@u~w�Op �E����h��p�����dT��'���rg:�l��ߛ;X9d,��^��e��[Kh�-`�9$~o������eR���E��+y���o7쀮��V�2d�u�?"8t�{jV������������	�2��IA2,�"�e���Y�.,��j�*�"(�]���<�ѓ�h�'�1�)E�Kk@+d��=��`�lm��� ��H�=�.�m��f�B:��jџ���~1m9(^�������C���L��?�����{�ӝ7)�*/���/�:$ч
�RSPZ�u��_���\���q1��^� 8]3/�3�-9�wٞ�)��	���Rl�t)� ��R��٣}%,'"���x��y%�KϠ[o��-	~W�SZ�����?�u��qY�g��ǌ�X�ڠ�g(θ�B�_Wtΰ��>5�2Ы�0sڏp*'�i�M� [E�ڜY'�\z�g�z�iR�2W?���#��ʔ���*-Tϗ������E�S���+&gy�8��H���.��+�`�B��^��.5�F�zY���
�Gun���#�k����1�%d�]d��Y������kFk��uB?�����c=��Q0`�z�n�4i@�M��^�D ��|s*�DcBu�ڏn�7r>x;O6�/Q��p���ξ� �0������& �O`�73=[@J�
d.r��i�|�;$�Z���A��Y����y!b���wb��HX9~B�U���o[�Y����6ª�Q���������fZ�:��BN��~{E"�������iH��FVdʥ��d���2��/���$z�������Z����.��*މ��� vW���P�j#�Tn�Ly�
ǘ7���{;)r�I�u[�; j��P9/A&��oK]�e|d���dRT&�y���-d£��'U,�٘e�7�h	s��O��S�@�|�W<uF�.tļ������,N��o��X��d�֩�L�6�G��hk�Y{}�c'TD�Η���f�]0�c�,��\ ��Ep����F�.�'4Żu?g��CK�s�(��(U!ac�3��i������-قf���2���̃�@���Y��W̰�ɂ��%s&�H�/�-�p1^%gO�'m �N�&�����#8�Qx.��jΒ����3���]DGO��zy����"%RJN�zp7��ԃ�9b���'-���ֵ�˸�N��.����P�4Jɗ�-R�K��l4J�-&3F��B�\�FFz�+�?̝U�0˖ا�~��7�Ix����tE-]��/���J���HN�.�MV"�GI��m���\�O����ċv�>��Dk�Q�k��J@��Q�sQZE3��������񪈪)T�S6���x�6Sû��P�$*�N�a���q�?׉�衞�s�*��)���g`D��:�ϵu`<�@�v����Zt�w��V6!�'EkN��g;�?xBɵ�	��x{�)��u(�}��5�����x;ߵ6��M��c��F������a�ZH-CW�$���TԱ�nN�,�Z�"}m14�.^����a�}V;"��}�<ZM�T��ät�|W=l���Î2�A; Λ�S�q���E|�|aǓ�	3ɹW��^,P��z�$���&4 �\K�c����L��9�m)�@i�}�G'Վ�"ߒ�=�h�K_�;�����(%0�r�������������k?������|��][vfD�o����/�o*ϊ�2� ��1_�Pu�A��F�~�S�������V��R�뿯ʎ(W�s��&w�E���E�3���BaN�h�Y���~�cS◓��h<8qn_���N�[ӡ��@��ސ�	�l�oI�\�n� �nm��?�G�t9ů��?�)�W �P��%^t������1�(��سw�Tq�pn�o$�*��=\�,2>�6֒o�ۻ(��������e��q�L	7�휲iM6�\O��2
;�T�C�I���hY���yIw��K�+��c����NX��֔O�y*�sG�,��!�:V����Nm��p�Tii��K�,�1���c�c�SCx��]H��Ϊ��aY%��'��t3܂��}��A�ₓ�^5�Ȯ6I>1x1`o��"�V�Xװ8�C� �NȎLf�\Mƴ\�o���/q'?@�u3٭p����S��/�{!A�/L�L�,�Î�*Ki���bi��|��;��U�ޱrOY㝅�����g*�^�
�gO@n�m� ����������
�^ƪ7���`,^	���<�0��%��m�C���0uڅIpA���r�V%g� M�"]��h��ϵ����|����z	(�Iy�?^�a�1h��^,�&�D�K�*.[I���\>\-Kz��A��h"�l,?��ΚD�Z~0�<�@eV�oo�����M��r5}Ǭ.�n0������.)�@�7��%y;����ӑqKH�����P|v�lO}L໶?|��%�<��<s��Ԑ�f����&=����u��q��I��n��ޱ�����8�#D"�2ʜ�6F�s��j��ˏ��&���)�M=��S9p�S� �/~��$w���7�Y�Ӓm�h�s� �@7��s��q߶9�w\��"qM���[����|����(/0���l(</-�zs��Z����T�a��`15fIM�7�O��i;�Ҍ�yq�a�m���S75���O�JO��F߂��������#,��ǖ�'5I�I��M��;�!�X7@R�n'���Z���Y5 b�`��B��S�3A��ۙ��̌1���е�{��)Oٗ���W�5�D|���b����!u$�O��o�dQ�u #>�c��^/���]�ɡ�-�k�!���������嗛���Ʉ���+��?Cg��jh����#�ޝ{���ͦ���K�D@�9��h�ˍ&��r)aG�j~��&�l�<Ӕ0��>������U%`I��ü���Rq�H��C���ws-��}q���q��Y�cv�P/�h�K�����C%���e�����Ld{���yS�	n�6���*z/�t	��t���Q�dP��j����gW=-��S�08��C�T}�m�q��]�`r8��${����E��H̟'%8�-�d�ۘ>.3����j�L�΀��5���U�,p�'%厵k���� ���p��_D��,�Eb~�KQ�H�G�r;�������m��O\
����^�&�Y�������8�dB<�6�6)�U8��Zy�>*�kl#�q�ý����*r�o��.L�aǾ�q��O�Oj��(�_���g�:���m<Vv���c�.snʔɴ����x�5�A��V�6ވ�Eq��(t&����/���X3��w2�����|��t���QGa�S+��۔���9�,�;i������WM�fV�ڌZ,G V6��:/#���1�٠鍰��e���� ��vr3���w"I�rL'e���Q���g��!��r}'@� H�苦j+����'פ�C����Z�.�y&̶l�!2]oQ߷ec����#/1�>!qb`"��	}��45��a��yu�� �d�r���o���B1�U#�� ~�I�Eq���"�KhF�	V{�s����C�s�=�����l<�}��XA�)ٜ4�/1ew��vp��k	QX�XG��VB�\JH�-��UZ��gHLO�U�̮��g��/��\�ui�i�l�cv���Wr�����!�@�s�l�)W`���؜�}S\����_$�,��z��d��09�-C�BS
�����vؓ�:��ئX
-ݑ�\"�١}�S���̒}��#`<����q�~vm�;5Ҧ�ćiM�-a��kIc��ۙ���>��yU�~��ۢɲǚs��:h�ms֕����y�T�1UQc�}v�߱�v�AE@ƞ���u�Σ���5�6��R�w���(m_q��KZ#��	s���yx�{ۻ"�� W-@欩eU��t��_�(��DY[�D�?�_��܎م��DD�U�Vf2��f�ۆ���TO��F���G��rI)��}�s��W��"�A��m�&_�s_��@&���Θ��nT����Wu��+.�]�L�]wOҳY���B��-.2*�(��4�z�L�)[���C r�"4{Y��t��f*$F����/����E�5����S����6������|��&
W�T^)���������/J]1�;��X89n!�����ۃ�P.!��j��r����m��nֳì��gqF߂;gN��w_�o�~eD�a�HP�t�ԯd����r>΃�!�k�u'q5���,���4�ϵM �	�f�G���~�V��y���#�i����L%\��D�)Xe�p�u�T�j�\T�G�Ǵ7`�N+���;��h�@r-�m����@�zq!'��0�X$�#�+�|n���eZ�2|^}�gDG��Y1ސ��>�0!�	Y�'̽'���4��b�$BL}u����R|�h������G�u�!��&c�z6�{,���MDۖx@�"��T* �\9�H��w�MI%�
$_zf��/�lH>^�B��L]@��ܽ�a��i�����s�$h_���zp
yҤ�����_�afz����\�fmf���.hkX�4~�71�>U���9�I@�:�*f.�a/W�I��7[d�/Թ�å�YQ�h�Ù��Qrr�_��S\��~�������wG�p���}�/8@T���! �/єt�ĝێ礡�Fb���f��1<�t%x�1YX�B8Hi�w�X۫η<�?T�v��;�#])4��|�������|j��-��� IrNy5R��H?����u}x)Q���㊆2n�SL�\j����\ٰRL\���Z�!��?r�kß.I���{����DH?<�!j��*"M�Yn�I�p]&�����_Rę���Vg�& '�@H� �8���nfyo���7��?�#��b�E�AK7ڑD0��~n���-�P�ʝA��֭И΄��f�"�T��5V���DtD�j�B1$�u�d��j��JQ��K�E��^T��kэ�m6 XG��f���՚��)����)w�<nN�E�!��D�T3n,�^ q�?AN���<*��=�T�}�.��x��Q�9���OY� d�r�Ω!�3���3��~��C�C�4��)�i�D��+`S��Q^�FWQ�5T��xk����	�F躲�)�ޟ����,9��[/��� �-�'h�����	4����*[�!�^``ˡ�6�a��6�֣��*�F*.���M��)5_�J���b�ٽǋ�<W��M����1ư� �{1��י���P�w�T���7e��]����+5�"�KXBҊf��J���?��SN�8��R��[N�GL	, ��l%m�Ko�v˦@YXɚ�7���rr��A�iy��@�h�2�N��[���j�&ޭQ�	 �#���:^A5��[�̆�~0�U��Ϸ�D�x*�	9���i'��s�%�]�IU�Wy�Դ��R���Xpu�yK@YD�%�g�E	̲$�*̿%;YZ�q�A��v���-	�G��}���Nh�\�MճR�ŃL��/N�!�n�\�á�����D��V��D.�>F��δ��g6�~���:-��&�=���/�[��$�2HRy�W��� �i����p�P�<�Z��g$B��C,��^k'�\/ �(-�oX���Dܣ�.�cK� L>��� �݁�Z��瘍#f�M�cf��B,��r�iJ
> GiJ��Q9����[R>��a���-�9H{�_��	#��Ol"��ž��;/���%��)�n;4<�01�'L,�n)�W�Pa��Z�r�/�C?#������-݌������o.��������7E�}6�E�B�D���ϫ���\��l �Q�!R�������x��Zcj�jf��"r�3�`Jj[�b�tr���4�7)���fEp�����+H	Ю��@ ��3��.��_��P�7Eݑ��ma(�ZA1��F�%�*�<�
.�㰴�Sw���X�V����ɠ9�b�F+��!Z�ͬ����7��xZ�wH�N�����Y����v�][jAY$�������f!9  �	tm#�x���l���$n)뱛���`4P�֝g����)N�j�T�~pk�6���;�8$y�w��# ���C8v�[%BDk�zS�	�v�6]1����f�������<�u)��H�0sL�G,�e�2��X�x	���fئ?�����$'7���{`��Κ�OZic�w�^_���r;�]J"���_Z	�O�����̒��\�����#3f��'4;��a�ß*�_�꾹���G`�<��ʺot�s�(�`�	����m�$�W�>����xp���Q�h2nf��K�\�xW+ai�2�)az�)C"W����ӫ�& ~�>�$���[������L�\�4M�o��<k������7f�)�?2����|�֖�d6��m�o!޿�����0��ܽ�ЋyK驲�Ez���� ���=f�H���2��P�吶HFn<}L���_���	n�9s�� X�+ϥ�kE��TV�ٝ��\q("�m�"o&��-�W���kb?�A�j��J$��j�0� petz������� �yY�#�90�
�1��0�Z�0U<h��b�C��n�f[�T��aK�Ghy�J�q|
�50����3�G��y��4,*�fS��j��=x��u�
�g�An�PvZ�Ȟ�F�O8��ə��@�Iz~��n��� M�ql�M���3l~y�5����X[2��>�iG$�m���&�BA�\���=��Z�Ca�Ը1$�q'(�3���K*߸�t#���.�|�]`L<]�ը�Y�jŢf��X� �vn'�k�P��q����u�������=X�,l&ǀ�cչ�����p�2��O�ĀY��l���9'kA�Rm����'U^��H%ӈ�̱Lƴ+�Q"?����K��]`e3��[6��^�9��6�������?j�탚��9X�������n�ǲj���C80�c�+K�?v^�G1TU[�(�JBǋ8�NQnVa�
`;�")���#�5f|^��ɼ�j���R3����2t��	R9_ĊM�x�3��LK�N�KB!Y@�q�k���$U�w��wl�8�\��4��5B�	A�}5@ju�$����'B��T��F�Mߏv�"~Ѷi�G8X�5+7FxB���h�Pߧe0R��z���slX�A��T��l�%�p�r4O��9�o���;b���td�{�o��5ο����r���/���v���Y���(���D����觊��[�|��"�3��@{�UE�U��17)���y���Ȃ�?|�.]cy��5�~�+#X[��Uߛ�L���ڦ]��kf����;��{ 6*m, �~Ld~��u����B#�˛��apZJSO:Ř�i���q��?�¢�|���<�PI�e�m}(��ey#��1z Z��5������:V�'Ɏ��N\��֠W�s�F�-�ʩ����n�"- l�\��+�}�@���n:A0��4�ym�2���se�}��MF�d��?J��{��Z9� �RX<��|;�c�0Lk���<����7 ��*�=r��ý�g�2�"8�Ng;�yؐ��r �Q5��(�=t�	ڛ�ph��|�C�eb^:<;�(Θ��L��@~3������&/Xp�$ʘ��y�Z-|5:�`.t�*o�;x1R��A��z���j��с���:���G�����0���cV�M�ot�&�Y-�l�&�(f���i��<�L���/)Y��/���oD<���됢����mKE��[���2����9�+�w~v���b�D]�;�6�~�TX��Ȉm�D�C�Jr�1k��d�vP�Z7��4k*Fu�\ymĲ��绥KZϻZ��{ƴ4�d�mQ"�&&���Ws껁�a�:xP�J89#��S���k���Q�G����Y��N�Q+)�[/62m�!�\8J�X@ҟW*��Vj$K��N8e�t�A�=6�cNLޘ�s~�/�<k��<�L��r��(�.��/���~���o�p����/
��3��@<��|W��B���%��N+V}<�rMZ�Ÿ�CXn�j�����*J��s�+�7�GR�DD�q�"7��hr�Z{=��ÚTŴ�'o�Y�^�Bv�x<�c<���`�%<��}�GQ����D��MA��6���d���NW�T-a�ؚ	���:�f�n�>�~�h���t�����W34��"��e;�'_l��:�:���)��pЍ����H|�V�XU��F�������Vo��\2p�z�Emc��k��w�n���
N�yE�\^���h�=�4��=.�_b�~q�-m]S~_ѐ<�c?��1�yJ{����'1����Q�v�g�w1!�!ܜ��Y's�Ȗq ��;�b�~�p�EL��[���fH�d"�m[ǻy;��IbG�_�̽ʗ9���2.w^�}k�*J��p���އk�a�]ٓ��M;�����k~!���Ԕ�|v�R�� 5�V^[U�{�/�~�ު�e���w``P�pNRsd��;k��J��¡���H?���e�=���l\�\�Z��9 �����ӒX��#�����f/�N8�d��2��y��/�Խ�m�f*I�g�*�Q�ͥ�9������ ���DT2r�4��t�����'0�� ��o������WC������u�((åE��e{a8�o7�2����9�һ��ܶ}��|>��9��s�K�#�ow��6d`�Yڞ��%� �zT�(N��[h)5zE� ��*���[��=�9�öu����!~�?�5TI���m��Ѩ��ظ�����
;�Q�"�ˣ�D�_���)o�S6��嫆�-���w˧q��x\��g�|�@�	�X�Lf/|��/����y�d�,Oko����N�,����·��f���1�Nb]��.�����{4^�f�]$�w�\�	;O$�ȶ8�q�k���|l
��v�v��ܵ�5هǷ��?os��������co�+�נ&��^$y�	�G��>r�ѥ��� M��Gb�2��#�G�AK��Q���1Z��}�˾I�*�Ț(�]��T���
�qG'��Ƹe�~�9�<�R�X�07�F�ȟm��p�9�d��M��J���_���g&�����Ƕ�������/r�<(��q<�ٻ��]����R���y��;2{���������]�=��U�,B��s�IU�j�`��B��̆���E߬��@�w�/�r���}y�x��B�
S^�г%��Ѓ"9ԝ���MDbJ��YÓ��T|&-��ߡ&HK�8�3�P�,8��1����=�c$�����n���Y���'ccQY�;�%	a���|T�������<T�3%�q��m
k
j�Y�?����Z$Fv1qO����d��9a��H7����
�:��+F���v>��T7��ў��p�J�>si�鶋����%���c�h�&����կ����-H�D���Ju�#�]���Mʕh[2��q���Le�yZ����;5�*��B�� �"�E��:t��]|*��)��ա`l톦�g�CWb[:8]�㶏=��J��։�@W�)
�!:nq1���eA��K�ǃp��?]��~5N9~w����)Wͫ���ӆ�u}����Ul��,8U��BW̕�ֽ�|#�;k�3FSf�h��_~���2{��>Sp��Q���k�c�ecfO�>�Ӛ�2�-wf��v�Ӱ���e�l3˧�AwdM�>�Y�p)�qr�ʠU��j�è�5nLr3�O����dW��܂'����L[�"���I�,a�
j��G[�>��6F7���Y��c���F�к 9�=�FcOOԽ3��o¶Y)`���O��a���)�x�f��Џ��� e�ѿ�D)dx-�!�3��+u�V5�]���㻔�aV�
TW���nmlP?���ס�C�E%�F��T��:�[��~�Y��$�� �b�U�N(��Mc��/��s���SF�X86��vm�Uq驹������{�B��f���))�ӳo�HU�*o�g�߷[��ne�N(P��¨�g؊�1:�l��h51 #�O�۝����H���u�{~�2�zR9��.�td�
���k���6̴��yzn'ı��{��5F�й aCP�xt���79I��z�)�{��Ƿ�7u&i&�!�D��I3�K���^Mڦ_6<��c�!�v*cPUT�C?�"�{bܩ��8u�O��퓹�r�����f���M¦�
~�v=��?����X�)�����?s����Iy43���?/���)-ΓÑ+CVx�n?���:����k0%�
L}Dv?���� �X��r��S{q7�R��I�}I��8���M��jT(��3��m88�ڑg�EdwX�h�=5��p������Q���S��g&������'@N��GГ�<<H^��O@�+��i�tJ�?��^Ģݽ
�?�~�T�̗Z��`Q'Á0s�>s@-|ŝ��&:�-�QB�_���5��B{��t�L(��1�(]ቈco�"�I�ZX�/�����i�T:⩤���vׇ���t�F5�d���+��jRY�X#��Wa���c2�gq��d�
Y՜���U�M�����`��O\��f��������v%�YP�b���eK�HuݮA�?�4N��<s�6���0D�Ɨb	�uX���)O�M�/=��[	8�u#�
�Yr�8����M�l��E1�dj�/u;w�ފ�Iax�N��\�:�0P�.�ʖ���t����WY�Ƙ�LP�5ȯ>6)qx�3���~4Z�{�5 �74esٖ`�v�0в LQ��}�����u�%����o%r�7	fܧRf�i��w����L�0�6�y��6ĩ�ֵ�$$�H~���KC�ˬD�d�E��B�A����o�1:_�C*7���BZ�,5U�?�n�������/�l�����"~_4��}sF��ԫ�j[�s�݋��(�L�&�^b}ҿw���(h<�����ibI_�:�!�6�@N��]U�7���@'����{uN>�ӄl�+Ñ��x6?�)�Q�T��f�d3�R9����/��s� =k+��D�:���.��<ȡ��8�19-�U���6�`�L���Ή���U��ρ����H�f�FҖ�3ab���W�P@ߌ���bLBu]��;��$s Eo��3(�V�/����L^�?�e�@7幻�B�8�O�5���t��ʌT��1��E��+����2�B�����U��c֕�P�e�
������щ�ܐ?���|��b��Hg#ޘ�@x ���P�("HAyܻ��`�� ���)�G��dC�)�;�m���s_� C��L����g�yR*5��,��b�,o��P>4�~��+�.Q��PK:�3�=rVfI��W��7��,�YC��E�Y�}��1��(�*e��<�wd�19�&[�~����D�
fx\f������S��: �{"/�_d�}r3g�^SR8?�ѦvF���r!Þ�����V��O�"�&�����Ur��U�kR=��G�_�f�;��q������ K�͈d�dD}*���í�=(߹�4��<]ǽɗ��M^n*E��O�����G��-h6�"@��)���H(�@`��έ��j(<�����/=�L�9�Ը�)�X�6��ߡ�Mq�� 猖w��)�|�Ӟ1�KJyQ��t�]�7�>�xlAGu� mͱ����pd1K������EHY�jy��yaX,��PcV8���P�(= �95�<��:b���K�B�מ�I	��h�EG����ţ;�0 ���B����П��� �ګ�4�z��o&��-�D�fa,��4���A�\-�������ib��B.�=D��R�h���a����L5���f�߁�;�q�m�(�泣�}��웳@o�鏓PD`)M��f��ϊ�/K�o����8�����}�;�!�0o O��abn��lH7UN��062ds5���9A�pId��"��Y��frX���mP_umqr
�<XZ���h]�#�F�!iLx*d��f .Ƒ�,��c�G�6�@��>P����yd�f����Zw���D����
�.�Vg��x;�Uaj[�j�Ī�!_B��H�_� f_ڋ�-���h'��U����\ e����1���q~�q�UV��f��;�`��2��UˑW1�
�E�P'�	 l.�JT��r�.���Ao�?�����~�E}�2��I�+�f��?Ɨ��r`�]��`���J�6dn������������ɸ��r�{��������d��U�ɩ@E�}�`:�h�=a{}g�7�������(7�F�
7��jEq� Ol�aE�͢�e�P��RWWk�(hi�����	�&�x�f)l������g��B�+���4O�]]�!����z���)�/�j��c����Vm������I�3�g�V���yZ����c2����|�?�Oŕ��8S��l��D��n|�R�� ũ$�ג�4'j7�������NoMC��M�N�|�\����M��GCnh"���M�c�-����?A��/��I]R�f��;���g+��T_��ښ��(��2��2F��˟�z[
r;o���.@����q�5>}M���v��< ��R~��0�u�8J����E���js���o���a�O��6#��d����[�;O���W�B�1�p�]�]�����|�xy)��4[A`%�-B$K��U�:P� �u�)��#�[�i���G�dIM��yHW�������P9�\Kw���y:X?�V|��,��P�a�%����`�>�Ŝ���R��5�_�,�x����r���6�Hd̫+	_��J%��y`GY^-~2~�AO5V���ִ�4���{j��q�~-)�����ʠ�k�I�L������w�!CSi�e�u�a G�S3e�0^޵�U��t��7��l��=�|él�X��z��Ѥ>�N�uN�6�yG9��3�%CQ�Gl�Ǿ[��)[��f�[�qV��&(53�m{��6��)���դ8�*�˱3C^i3�5
uf��RMܗ�j�4DS��?�7��|ݙ*��u#���o1Z���(��Nd�ȯØbC�a�����"��T�58H_T"_��%�;�z[7����ݡ|rD6��a����2o���/@����xC�_�P��{���Ĺ�s�#N��0�6���Ƌ-.�dg��4˯.�J��P�?���Q��`��Q�ۦ�R�
TQ�ε�8��L	H�*�Nwz�#��r���=Āb	0t�盰�=aBU���5>�7��g����'��0)�<
�b���8yv�$���Ȅu� ټ4�8�R*'%��H�b��rVP㧊K_�Mv���M��+`��Og��9�x8�w'��G\��` .���.�j�6ˢ��|���q���;�"�/��&iW���ӕ2@�F{��R:�@���q3�3��AFHA��E���
Ԙ1)�0A��\%���^u<;U��-���M3�*Qg��ɘ��M,U��Կ�tν�^�彤j��|�.Z%+0eS6Oa�|݋�V3\LSҷS�c����Q��5�R����lg2�T5!v��7���G�A���^��P^*MLKFM�B�J��:��J�ω����;T���l�g�/�0mgw��D��-�����Oւ����^�F���\˒u^��Ы��1�G��b�|L��LHDI_��݁߰��{kn��R������y�};���Nu����zR�3IV!p6��C���m����:X)}T��k�*�eT��\��XE�=��t��}ju�9���*r�A�E��V��8�2z3:Y�tj��ٺ����c���ޝ����ȤjUR��E�Q�傈6�^m�7j_D�������Y�Â�����]&�{R�b1�oubl1#��3k��,�s���=1�`��~k�@8!��ƅRX�Oul]<j|����\��$�-9ht
ۂ(��T�Pb�lz��gn�!��T�3��@zx��I�WsG�Y�,D9�UUPu %>1�F/�L8^�=z��T{�bWS�4��@a�t�A�xQ�O���r�\al�x�/ʩv�`j]j=�S?��:��������K4�_�����Le���8Èb�B[��&�p>E����ԋXGJt�
8�J�h�^ˉ<��� ���hG�d�O���U�N�� 4��2%���>c�.X������D��֣�9��T#"y��7e��3|�H%#���.�i'8MSi=�*v(Y��w�K�$h��:����$�RrKؿ�vP}l&^�*�R�_N4���,r(��(�H��Ӂ9
9�3*��d|�R���g~-��4u�k��a:֭�]b��s���p���W�8����E>lSõ���ޭ[�?�CL �'�?�����_�1��K�Șuζ�j1�4�Ec��9��]ުrX�B�?-5�Ӓn(�5�3����R ����8�;�y6L� ;N���T�T����&�䵲�&)»��|��:ޤ�N�l�2K�	�ڙ=��b*�ke�j�1��)����b�0�I�l���k!��������M� zS�2�9O:"V�IzRG-�G���X䚓�¦�[�Z��5�l�ptc`�옳ܿԕϥΌYÜY��b0�&66g�R�y�Y�?�m�A_�4piޔ$Yu�¤�z*���2��BU
�v��sܽ�M�E����s��qs��Ҡ(�/���sG_K�`=�����My�xU&�P�Eî�^��b�8;8��HF���g�\��lu��18e�W$&b �5�)˄��N�|\T/�5?M���ɰ�{�x�M�>\0�ȉ�!X�8����=�LQ�3Z�p�-YQ��u��j��;��2�����	jkw���r�����b����7��l��ߑxή#�vy�,~��5<�G��K��N�<(]<���耉'���T[Ry��\qN̈�W�~Pj~��YP߀�s���Q��.��C��-޷d���0����F,g�� ���� I�jMf������} �d`+�8���D�W8�!Q-�9
ۚ��2+_v�3g� �he���s��A����lhA�]�>W�#E[ak���3��8��l�G�
!���������:!.=�hk��涼:�-��0A�Gr���Q�p)8�|�Ջ��т���Szs�l�\1�޷&|�Vgu��!��!��ں
'��ԲE�i�����Xi[��	���ȇ���b�SF�d�׸�%�����'}��ғ�3]�:�c�+�H��΄P� e��zw����̓o�~�u�~���u�*ͨ�q����[F��M�&C=G�(�ˣ�03�O�Z�&�|r�q��bn=��I�?t���V}wӭ+�^���sԔF\+C?��<�
%yFчyg����"�� ��ec�n,����]������S"��[�B�������CWҔg	#��Υ�E��*�j?��J�w�k�Ai�;8���ג��3���f�qq\��V��� ���
�l۩.~���Ql���<�����bD�(�CK��W���g
��2�ad�m#21}%�*�0Ii8��$5�����1�0[$^gW��N=o�g�n>{�cb�p	h��t�?6: s�j�(��o�k��tCF��]>Qlt�{@>����_���9=����J�ϮLe�I���Ta!���T�u�QEL��(��!}�`?y�j�A}�YF�����Ia:��7�auv,�$�	�3��ndxg��i�*!g� 𧒁i��PY�P��?V'�<{o����r�r,}5��bk���P��x��k��.)������>��F�!q��_o���>�XN�����$:�T� � �J �^���˗H���{�r��7B���ݖ<��Pۀ�8ޕ��F	��坻6��%�*�������6S6��%x��<oa(s�utD4l���wp��)!l�5&����X����C���:�6��L�������qr�n���������m��
W���W{B��Z�a�{-���L�P�46��/��]f�3g�ʡ5pJ�.���s�f�j�<��}���@.��@,�_��C7��Z<A	��م���U��٬�ƥ|�<gջ���=�Ahx�HF5V,�.�\�u�0�+�2���=G�8Ԅ3ŝ���ۀo����
��J.SB�l����#).0� �O��>ϡS-���A��<Pp$�@���� ��)f�7E��NGNF�GM��<^Hi�'T��\Ra�^]_<�bl�V���>vP˥+��@�;Δ��Pc�:����r�+F;����g1s���wD�<��Tܾۊ$�����}Q����ƙ���՘�D{��;�)t����4�8��"Z����?�U6-��{�=�vi�}<��p�v�=�� ��&�_N1z�Z��]nU�f"K߄{Rk��)������1�8O VPC�<�w/�HH��:��`@f�
�i�f����n��ྫྷ���=0�]�{eK>|��O�M���_��ر��G^�����TD���{�ee\����r��=<��c���v���e�A] @̰���w�3�ZJ�+sn�@+ǼVK�C�� v�r���J
��n�G�ng`�|`B����C�a@��r��TM�T&Ź�m]��r�jhw<!&>��Wt%q"m{�2l��4V��D��1�z��~p|�0�`��;����kB~x����l�/>wً±0��3��z���"�޸�_e��r{c�8r��v��Ro:us2��2D�	�"w� =$�֌L���5�0_P�y�VH�N���H�_��Wʱ�L�����xiuJF�6����d[}%�J®�t����-4A���U��/� ~�`��(��Q���o7�|�@�L��=F�m�����Gr=����߯
O���aL�	f�L��^YZ��9 ���u�h�&�R��n�ܲ�3�]�g��<� �E��+L�J:�Ό�t�]�Ĩ�4�Oy��p/�����,�p�G��Ą4 ͋/�aSRx�$H���f7�E�ʧ�A!!93S��nNZ��0�v�z�k��.>�u9w�e,�����5��8ذf�C��>�W�W�Εb?����4fס}I6��Ȣ�$�lz��{4_z�.T���k�)]�)b)�0yk���KX��:E��Ħ��J����U	./��>%�M-�ir/���^s>yg2�����������f�N��:T-$�0Z8��-���3�<҆�,��0���6�.1M�?�̘"1J���p����#b�-�����.�V-�V�)ԁ�գ픲;'1�"��w�_T.�������
:����͛O��n���;��6x�uiw����[=�ۮY���Z�������]��M� �]?��dBGe�v��y�`֫��>���x��4)>Ӳb���q�͐��)�X�Od�>�T����N��ׯ�W�OW����y�����Й�bp+����O�!�͂1Hm��bVY7ס�u�ex�I��b_`1_�K7��CoJ�!b�-5˃�<�����"���up@<5~�����u�i�Gڂ4��=�h��~�,�h&(h�T�B;J�����w���Lx����?��'�c���������2���٦��A[m*�B6�G!@��-{尳j��V+�����mB�1�"�	zߑ${��6�����Nh���{�M��Ң��``���E�jqJL����2FĊ���g����@�t"</�^�{��}Ò��|�<���N���U�.a�����GtA���̱�{zaQJ
����T����c|���B1wq���6x�'��[�ȏʱ�K_#�G���2��b0�jI�]$�~"M�j<h�%��J���xY�ey_��^�n���R��j�1���o�8�XrC�2�Ò���,�������!*�}D���v�{h+j ��ٌ^���>�J*��_�����bp3o�$��`����w��Җ�/B�iM�xZ��
�>MK���5���DT�PH�n��tE�B?��K��VCo�#�-�*��2^8��Wc0 �S޾P�b���YTg��-��|�G�����
��&B����#nt�ڎ���ӣTԵ���u �`�<B:_� ��'
,&:ˣG��_��M2qL���[�]1����E/��"�o�j��2/���o~Ln��dW"Ud �{�~:�zv�$M�^�l��gW�A4?������{<�Kg�_Ugw�f�\ŏS�֔�ӝ�߄����p��y�5]$\|���=�KD_g�}홚�"�йG��s)��ah6�č�kW���"�/NP�
�V�k�e^�;�Y�}���sI�d�9n�brL���?��ˋ3�d�����:y2'����B��ii��,�f����_�Q��%�j���C,x9ES�a�b$�J�����3^�~5<�Ze��H�i�H	t��u���Ա����"X�I[�&_���4�A$�;)�3��c8@g>
��x�4o�Jr��ñ7��\2P�J5�g�?��6���]a���SΎ�͘ �Y O%-�U��F8�ċx��*��H-P?7Lø�[�Ty �`��]Ol��(�!`�/��E��F��X�.  +"��oX����+�?�j�(B|�R��I����M��BU��8$���VD;K�6h�,L�f�>���I2a�L��ᵟ�ژ�m�;�:�!��R��N�����q��pbm�Zj�	E����L8W��E�c���k����)R4% �!>��=	�9���$e#�ۣ�ót&6�|�)_�k�r�d��>U��<�����������[�:�>�BT�C.�8�7`Ų�8�$�� k��"���H�����Tמ� ʠ�>�m���M�<�%�ja��lΕ��|�Ζ4��F�����N�=�@
_��ң��5_�4��LF�+r�{�ue$����!n��zlV�N�E��B�d�)��?��s�����嵿a����u�0�E�������UUW���o���/� �-��t9��`Fu�b���!pn�QlN*�����X=����n�b�z�x�mg��+Q������TG��׉�t�G�ml�3���JF>���ݟߤ�
��P>��>�N���E˲�W�c��3�*=Vqc�@��b+�����<�7H��;b.�
�P��`c�x��!���3�f����^��(�\]��$FTg�5��j������!�2��j0�e�:����[w�WRg�����X����m&<Nb_e���;��{pi��k%ayzZ �"W��[
�$��w>\�E�w:E��Y�UnlR�X����<����Y����Np@%�����	��#�Z�B�Rx�vr�q+̨�����g�y����{o�V�҄�oE���DAso�I>"P1<��e�Ջ��Ln;C{^�	�.�y�&�iU�8t�>�L�y·O򟤶{y�=6��1��?�Wo{Bɣ�E�
�=F/CD]����D�]�@��hRmn�.�ڷ墹�Du^Gy�=���u�'�$�	���-V�tD��3�Y,EFT��V�RF���3m_�u�c��l��Y\+p���h�Aqu�Q�n�Z�j=A�l`{Uml���QlϨ�� V{���<*��;�ik��L���f�<��^y�v������<�O�9m��8������q�~��V��i.Aƣ��`&3b��9Vk�l'J?���rd�N3H� OA�(7Z����!$�����F���Lh�n��U���߱8�͙��?Wv�����.YW+��ت��ZexD�txz"�B|�9������52�����`b�HO�ӝ���36���n�8�%G-IÅ1��/�}�����R��˩x~�w,I}��ބ�$��;����%�QP^4n̂�΂yG��$�n ?���P?z� �5������ǫټ�d]P�I�Q��di-ɡK�\�yYE��D%���pH�p�k��]�AF,�z�IV)z�gcO[�≌��xm�����H2t�Z�L�*���UQ�5��tq�y!9�X<S`�T�+c�*�vw��R7����L,;0������'�����KR�Oԟ�IqЯAMy&��Q���)m5�|�OD�a�И���.�vu@�p�E�P�4K�vȓz3h�~&��a������CX�BM�ԍ�	�Ľ@|^�dʽEuG��;/�����;=T������F�������s"H&��.z�jwσ D�#n���3�	��Y�g�G��-͗Yp�z�q9���+-�IQ9��>��'E�[a6n4�U��ˌO�$$T��%��,:f"�C9X��e����lm!�	���!��L�8V"��45�O�b?+n�����Aa�v��$˙��#|� u��3�M���,D�~�V]?�6����l�C���A"u��È���-���������h�V�/Qmjlg1$���ocZ�q`t����ە����7����N~�D�
��ų�$�� ����mw��F7ܨR����@�:��Ѡ����ri5��U��gI~*%��'�(T.��T�Y�S7\������{{��,���>0�ਤ`���:�m��C��A�O�����Y	�'�<�T{:t�r�e�fj6D}��S����6w�.&�H�vВ9�`�-�,�.��
��m��pMNn�f�U�s�87`���g��i���o�1��jm=x��lV\���)��f�ӣ]�����@�3�K�� }W����𫾈'�p�<�7)G�O�v��?��M�
`�@,�����:�����%���B��k�l�x(�����}���{�:��6��h&{��-�qx�*��V��ܗݮ ���w�,�'�� l��c���[�)Q�'����Z0}̪c�"��Eq G�|�`AZ��TLp���z��N����a�^(��O�n��6<Xz@�ꃁ������p,�������@��ϸ�}z_�����c\�
�F��/m�0,#8��g�h��w G4̋��gm�t��u��(��1k.@��H����hvr���޽�X�'���e�Naz�y�l<�eDT`�:��䲶&#�D���C��s�es�ǫi�����;�A�~��ꪨJ�Y�9��ϱ#I�|�qVw�u�h�xݖ$�0�nn�
!3�ǫ�Ӊ����ǹ� d����%�ҹ.>42�9��8��Q�q�x�2��� Û?wq�V���Q������{�[�S�3m�eu����lC�K��d��4��C��L`��	S`L��p��=�{�+���5��$[���gX�cG����Z.0Q9B�
O��r�}$2��� ���)�� 	n�j͐�>Ne�y�{�'���(D��T�^F���՞+}�<�*���H�F���y��b��kz�=�,�j��<����e_f!�]�,7?��f��\QG*t��o9[����e�F<��M�Amm�?~�$���XbUl�C=H���Yi����������z,���{����K:%v�Ы7�V���4퉠� Y�>#�Չ`m�)xЇf��Ǭ�x�����3�!B`Z��B/܌�fA�E��`�'!9eQ��%ϋp�-��d�2�v�V�c��U�w�e{Iux�)i�-om� ]d�`�ţ���� �}%��=�D��Ŧ�^�3,ϲs�QAU��+Ҭ4t��;q/��-'�x�|/(���\�ϥz�i�mp�@��5����{!����	��R>	ODݴ,a�+���jH�;��.�\�1eR���eJ�l�N�0�K����h��K̥S��ȵ��<7��U�j7èp�`"Mܐ��D}��q�&3���xP�󡣖�{ƃ�SL�N��.�XE�cG.�����&�!|l��� �|� �EAZeb"Ɔ�"oG�*?�MƮx��*eY}����b���q��.��} ��abӀ�]�e5��I2��.ϰJЃ���5T�@���$�K�x�c7�Y�?�rK����@K�%������E�?S�I��QՉ��)Q��S��c��j�eJ�.+k�8��+�T������ �,a�-TG���i��(8T��&'���Ѓ҂aHY�l��`W�?߉��C�H�e ��2��#N�g[�6�}���+{����#�Ln��%<X��2rH	L��?E����b�v�Hn����)�BH��^U=�3���T�,��~]܎PUƸ� ^�q���`��^�a�Dn�'����ۄi�񱴰R��t'v��;�*