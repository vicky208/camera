��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V�}��>��P�|_>ߏ�uћ�tZkt���&����hqI��^�~��=�@ =�B���d�1��|¾;��>��\:�O �R���ګl]�l�H�.4���|�M�����]?*\{���q`R{��R4Y�	J��>�<�����8m^��_@�L2�VEҲ.�3��JOԶiTn�*�H��\+��`2w���@�v${�w�~��ۉ�J���yjӪ�����
�`�B�G���ZX���xl@�(9$=E�ٴ/��ڼ����<C��.)�%���Lz�xzE3�"?*��Fj�d����=d
��
��������)�D/Bo=m)V�8��o-���n�{�#�NV�R,����Z�FHw��!��-��1���4E6�l�l-��5F��@�<2�.�h7=�����pi�q�E��Љ9�o�����3_X>�>r./_�1iAiI'ؖؼ-�Hg_�^{�p��v�k8U�ӮJA=���C#r�f���I,Hqi�5�'t#��i���27�4}��)�{��w����p�t�ЯMn;�.��"�������2� F8(�9���@fÊ?�;�:��S�� ��]�
a�� ��+�xB�
�N�Mm�3�-�J��p�`2�ӝ���)8��z ��j�|}�f`�(�C��+����r!���7�p,)�� M�ܗ��|5�g= ��.��Y�1�f~o��!H�0��ǽ7��pf�ugEI� /�oD�?V��}R.���$������^�s��>�^S�_*��	M�țZRO	�������!����Ouk���1ޏ=�W�7�R��:k08]&�6�j�����a�q�$@12cw�V��N/� !�N�E����ޠ���dy�/��ܜ�h��mʷQŧ�N,�U�������T�2�~֠��w�t�1�Te��-.�i	"(���W����b����n���Zt$f�襂��ዮ�d���/:���+��9Ŝ���(o�~/�\��V�H� �ɵe4�|r\Gח�"����^�Ϸ.,)	��c�l�?�r'���?��5�4ʘ�pU͝�� �q��N�$����wX�&������� �b%O�|�-���ܐ�Q1;~�^�X�&_A, y%`N�k0��c��5S�!S�i}]	��q�X�)Cщn �i��}��F���U[S��_�Ӈ� ~�\D��φyn���:��i���JT� �J�w�I��8���Rz�(��2!�����4 ���r�B,�Tvk����SY���cg'��Y1L���!1feؾm�q�tz������I�u��2L�ń+s����RK�S? ��6�=��c��x��Te�BH�%@�W�wx�x�^
��D߮_��j���^�;1rYEf��	�:���/��n���q�K���0�%l>!R���Q!���ca%����&b�+�qޟJ}���;)��@]�k^`� 7���TMcl2"�����)oH�A���;P�"q�2��|��ekxu�/�h�Zz���3�US]�}�C���uBLc�u���w��s�Gd_؂�ӕ��nf��_���"�)�K�-wC�t8����J���k[8E]åh�G�̍lwM�Ē��K�$zT7dއЖ�-�GpS��	���n��g�S�g��=�B�U�U+�k,����$��"حyȦ��
�qp��u\�#�qY�!�������Ky�ha�Z��	�ZH�aA��)W���m'@̌[v��(Ö&�)�����N��ysX�e@.E{�V�G�:��i��^��f����q���p�(;P	��f�0�Ir�
�L���f	�ג�;)�&�u$8��?�j�#"�[����M�~��D�w>���,�t�B�'�>0�C:�v����b����)�i��'jT{��ꋺ᷶.y\�*RMK~|fu3t�@i�*N��/y:?��䔨=�go��z�"��b&���ZJ/��Z�p�7@����'*C���'�0O�G]�}|b4�����ʃ��[{��lJ��i����ML����@ƥ��B�iIb%Ɯ�CziN�r,��:-��.�h�x�a���[k�1C�i�	��gk��g�BE�dr�����~"<N\8I��X�+p}
S���ޖ]e�^���N'V=���"&���!��׆�S�QCq<R	�UzF6����[y�EY*���f�Ű����/��v1�}��z��0��)�'���]����:�ɮ�W
s)���>:��t0^��׭�_��E��N�ܑ����BoQ��d��p�����h1�0�P�o��\ҭ�D�Bz൰g���߅� ���:��]��ꍖ�[�U"
(��*��L%���c,m��l� ������S �A=�f�e���զ$Š�����f>M����](�U2�~]s����"`��2�}ͻ�e�	*&zR8�V�@>�X����EUΟ�^0� �Iao�˕���Ϲv�����K���2�5d%�&x�)�I�59��l!@	�]�#g�5���W
	���	D#���q� A�xqє��s��D�}4L��zt���L�ʡbH�E[e������&�����L�
K�����(h��G��_��d�6��k����߭�Y|23n {˾V�զ��p�򮽔��h��?4Fn�%���X���桇qĤ��d��3=�X�s�Q�W�C��v�	�9L�ְ~�풿�}r�;��.���l�B�q(�n�hA!��ڐ�KC���t��'���-��X*&�eHɏ�ጹ�+	7�Y�~˪��A�	�v��{�ye������&:	ظR`j;F�z�z�F�a`T�������
c��|J�d��Me#Njæh>��f�ot`��z�tI�=}��؝.�j���^/u<��I���Kch<���.8�͙�톧��Y�sӬ�mtQ?����F��fN�#�!MD����}�)+7�5?��u��]��=����;C&���O�I�y%�ӟ�gO7��B�D>���w7�1�q�O��}IΕ�r+iVpĳ
�{��G�����2�_��xf��À�X�>n'�H�-�n^���$�B��J��I�-�{O�C*tDW�Ax��'��w�_����L@�/Ȭ�35+��:�N)���8u�\��!����b������Qi�?8�Ɂ)TV/W*O�?�/��踣O]��Z�٨�l�����PCX|i�3�v<�$b!�l���Um<���6�}g��+��3G�R�+����:��@jD?��a���FYI�
:K��2>���y�]�]��@�R��X�c�a���x���ݔ&nY棱��da����r���(� ei�=gO��G���CA,('+�»�ɗ-�9U_��,��^��裡������٘.�:ZE6&�5���������6WH��NiXM@+���Ahj3��΋�
����<�nv	�����I�p�/�>�)Rm#��p��!��U'kgf�c�HPfÝ+�Y��Ì��~q���]��ƔR_p���!�/eN�	���<9}�X�u�Im��F��̭�`_m��J��َ�wɚ�2�@�����wÓ|K�U�b����?V;�5W�9����2�=>�����uF�������#�'�*n�|�Jk�)̀��W�	c�=xԈ�<���|�[?py�1�$�G2]�o�)�b���r⒊_2MD�o8�m��,�0�"p)Y�m7_�S=P�(.�N4��3s��ogwm�;����yh�i,"�.�K�yS�@l���N2������ϡ��7�$w:��CÜ�0 �69�s��F�
�~��������	�ӍW?T�ކ ����!����$l%�vK\�ƥ/���~9��ڐ�$�q�n����FI��X�)�����+�u-$Te?�O�h���N!(PװY=.
	�����5Ϛ��7��EJ�X�k�+h�?|��/6�F\GW�pD�H��_�c��Ж4y���z�m�8����/����qO7oF����|��?H"�����#�z~���p��r��a�jAqC"��X�"�
t8_�9QYqQ��:A%�m=�?���݉ ����>Q8ܠu8rͤa�,*
�P��hج
�ۤ4!�:h��6��ۅ�Y�H�C��)�k��k�^F�=�ۉ=X�el�����j�h�s5F����/p���<a�zF�����압{{�UvjY�9���y�-�L裰՛�{�"�B8��� ?cs6��=5��)�";yן	���>I��zM����7k0|�������D�UD���W'�Tץ������-���D�1���/|��Ήh���2���!��������.�|
ٔHzM������q� �V!�t�DU��{�8�J��=W%*�A�y}	\�D���Ի���f2Ev!Y��H��k�e-e)�J�?���*Ӕ2��� >��9�!Q����>�3s��6�wf��F�꧰9`�q��2����a��\�	�?�2�l������1��ie��Ɛl��L�aq���J˞l!�R�'�$@{����z��S'dnX����ǣ�{��t*F�0�(s�6]�����*��\D%��~N�ǿ����O/��!~,=�)h+v� �Ƹ��?�-Y�V�P�߅�?z%�DV��H<��悅|����>�邔�NB�-H"�Y�iC�;b&�Y��m<�u�8CΕ��C��:��h��� i�S@���C��ڸ�\�K�X
@L�������ᶗa��r��X��&�gϭ/����%����Ih��댞��^lh�	�x�	̓�~���v��v�Id���aT&@���H�������c;f�<&�O!4���u ~�A�H%~��~qH�ܥ��+R .tۘ�����&�8=�ЙqAW���*�l��DqZG��}�� ֨��1�n+�i�l	�i�=U���Z�]�'�\Z������+���y�vn!�\t@��"
/�P~�:C�4?���q�Ph�yk�d�W_���M+�n�&�b�#��|��9����C-�����O��g�e��3�����M��;���56#7�'Xlp#R���r	J+������>��p&��F�����捪D���F�:όo�F�Oڧ�1Q.����tu��������Y�A�:��]7_���D+��[�7���OX������.�J��pK"��?��ARa�Z�W��\ ���\�{)h-�4�F�8����3�-�	o��6b�)&,����~�ח��t9oCkҞ}j�}Ot�Z\�����":�bQ��Pg���d_��q�-V�i����4ګt	wb� ��B;`���O����;���.��y�^R̞Wj��*��,]ԛ?{Rh�bL�!��j*xH���������� F�V�(�^��i�Z'N{N������R�\�*���bN�Am���Eܓ�e��p��vi�'U���٣���n(U�8M�q1�"���vZ�5N]���M����V����&������4��/h`��*`%`��� ��<���WXT�0���*u�N�¹���X���#7�y��Y�,+){8���W�������쵐��l:Cͧ�~6X�Fj�o�^r���"��B5*'}Ϡu_X �+Zp�GB�~�G�vuӟ49?{-��؍�%ļG���Cn���ү�oA��@ZMX�tIP���X��d	Ӆ�jI�$�����9����q@'>��<��#Q(�v�X"v�Ua�I��ݫc��$5^�pnʣ�}�З���'�s�㋙M��HN#:�%a��;W:�gs�B�#3Go����y�ѧ�Հ=O�0kcZĖ�sT�R�~Hf_�h"�'����O�k�z��j	p�<-fC��p[���x5�dk�uR{/��� r	���2���x��g4���H��7(�r���2#[!o�S@�� D|�Z_l��6���!y�.	p��1*[?��r�^J��*�_�󞤴���?OS#��g)%$��'�#;��(��q[���Ï��J_CkxL�q\�퓈i�Lb����C��wsޗ��
��"�G]��,��C�Ti�:9��~G��W��|�(/-�=�s;����yL;�/Fvw~ir��P��}�񕾦or�Ĵc��?Ϻ�F�$	Da0��?p��ǘ�N4�&��A���9,:Wp5jI��R ��9��<߈-WxX��EDԴ5')����@�����[>ø��d�������f[C+��ُ$K7կ�9b��U��?¶�t��(�4���9܅h_q��P��ܟ��r)7���ܺ��1.�!drᅉ�3�ş2�l[gR��=3��ϯ"�&�.a��J���KH��z��y�Ůi���U�H���4c��
$/�B��p�,��m���M5ҕa����e�<���Ҷ-��	+A����Q�cq�g��?�̙Q����;]��Z@60*U�_���@�ä����s���X��2�fY��	Պi %B��*�f#m�<�n"_~������7�7�� (�٩0��V��H�72ݓ y��=�j��3�N�tr�k��s�b����_�1�g�x�9�̓0Όk�y-w�\_��{��sď���N�ꈐ����|��{C��Y)��L��'V���/x��)�vo<���,��3�W�F�Ĕ��,������V��
���4���w�5��J*]�D@�/a֓"�C �HΎ�7�&�3��pd i�����{���h�z����K��b�
!,<�|ϥ��O,kƸVpH�e�cmq2���`���߿���SYhE0#����\L�3V9�e�=�+�ځ�^������6E�b:��R46O)l��(\3n�i�Jq����HCm����`�-�{��v�E��k��[�\��$��Gr�6�̪�C�"n��bD�������G��(.�'\��M,���%�=��6��݀w3|�"�^0o��<���w��"{?6A��c�J���R�\U�2f�7S�%���\g 3#y	� �G��� �3�=���B�U$�	R����1��J� `��˭�Gį�JÝ� �Om]��%�W=���^ź�qK_���3/jER�J\|4�mf�(�T-��W�K}�~�
C��0�����Ⱦ�<\���a�a;�|ۋ��?�q�5�Jw���ooM�%f(��=��pdFj�[�mڋ��!�Ȱ!$����J�A{�"\������\���Y��G�OM�˅[��Ql�:^M�ƹ��k8���p��g�T�m�xR�=���R�YҶ ;��CJ��E3��C����2i��t!G:��m��x�|%������m�@�x-��n=�tV~�g)�L���*�jA�xý��@�ya�L�C���^�\�RD=6�c�,)�:�I��>2��*|gN�Q7|��[�VX9 �m�;ȁ���-��R���ʨ@��I�c+�mF���	`�����*a�������;�Aŷ�^�jNq��aN���7�衞�{��]H��}�Ӡ>�&�W,� TW=��S�T�e������$����{�n����u�FU�J�r��sPϮPߍ�+cB65.h�-�~V�(J�"����D������K�W �����~v-�%�!F3�����"�%ٽ�b$Cl_��K�V.1ޢ�g~v�;��Ԧ㢺�P���&�nR�I}R�bO�Lɠ�p/6e�Q�%��W4�A�����Ҵ�T0r8������,Rb/�kp����n�{�go� ��E ��S��Y%ig�"*"xv󃑦�u�� z�&�Q ��t�m7�E�� �D�������t|��߇�T���"{ W��v��"���;f�8�P��I���-�xz7W�i7��w���6��i�q� %+�˙���xG�����ȱ�}`/��$�T=5�2�.h���7�Y���l��/����A���W�j�
8�Kg)�$�d9�I	�^ށ��Or�ɇa��t��R�N2��b�����/)�8����viu	:�5��q�9���@ ��V�q�V$�Bfk86O�*M/|�˭���]���<�M�%Fp]���s�!s���I����.n�`yoc���*�>^4� >
����e�!�ۆ�����ȩC���d#�7�-U3�[��c7�xͮ�$���-,zzS"&y���1VZ�*��L�b3Ձw~���ZM���]I�Q{�CR����{�bb��_k��-�\]Q�<�I�#ܒAf��_Zɕ��x��Pm�荕l���.k�3Y���s������b&���z�j�ۅ��� ?����΅�;22���@� ]@|�goƇL2r'�����9�w[�r�����cr���Z���[�ǂ4s�����ڠG�+Ol�SR!�
�'����ܸo�:�X{� 򪵥ݍT	�@
�is���j"B���qK'3�p����
"Cr