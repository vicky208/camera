��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�GN�Џ	�Ue�y� �o�naD�1>�z����Ȩ���x��<�Z��3B�,�*���i8!☞����X��eyؼ�U�$�Q�N9�Þ�tm�]t6���j�+�s@*�	VP�{��@���A�p�M�i�z�B����ˆ����+�${�Ħ*s_�cB��Z���C G����,M3Z�/��$0)@����j?t��9�0bHm��T�ƾF���X"*��n{/��Y���'t��|^zn�U���Y}\2]UXsqe�K;�"�Q�F�<E^[v�;��6�g��&5��(`�>.l���f�Q@<&J�AwG���P26m��2�GN��Ǌ3�9m�5B ȉ��?�����Γ����j'���"��I������6�TH�f`⬶!��Iצ�D�g<�����"r���.�P��4��Sք�J���r*�2��7�/y�HB�����������=o$�h!ۣ�#C�XR*���B�z�Χ,2� 8O��\Tܠ�9�0�b��P�ɩI:1���a����,�Z�� �����GȬ�O67��D�3��|�Z�޵�� �9��i�%}Yba���7��8��x���F�207ދ�����x><C,��7y����ۢ1�RF+2��VVS����/}b I�Ȯb7*b�\�(Ҏâ�*�/\�֠;�w�}_J�M�:�!l�a�LՂ�~^��AG��~����a@0�+_	MI��39	�7���,jd�L1��_��W��=f�����X=@?Zbn��6P���U�L����I�Z?��d�|K���	��t���1n`���WMD��_�#�G�"Ԕ�IIy5���Բ8��c`��uE�*�"ܧq$����<9�cf����u̔í�'$�)�"�V� =�Ӷ�&�*���ڗ��Zc�K��g]�d��Ԃ��{�a����}وrl$�o��!f�g��o���ME{P�,cAr�xtSi��nS��˻�d����-CA�L$X�}^Y�Z���rΙN��
b,{<&�Bǩ�Gh���0��u���eYy�>�,�el�
��+�7�R5^�!�q� H�~�������䏤RU�������������P�ua�Ŀl�Y�Ć���EF6m���t�-�R�6��-v=�RgJ�,��E��}��3K|��!���1s��+/M�q��:�<�C��Gύ�Ei�ң'�� �{x�E��9Ww����V���aR���3gz+v�E7�l�ǟ�d	�M�wX��"jM&P�{�o4��^mb��è����7�/9S�%��/����k�ͽ��Ym��0ٺ�����;�%���5z��"%�����$$��e������i�u��#�4��6����p��0[�%�1���[��#p����-��b�O/q� V�_��\��b�>f
�QK�_�{�?$g(�7�xg �k����5R�<ȸ�S���[��uoh#����|M����t���Ͱ�������J�!!��㉤;��Y��Q���)�Ʈ�ۉЋE>\Yp	h��[��'�ً^���>�kǭ-�Y*d�t���~�\���\��9��،ў-"K�Z50Q�ک ũV�QW.u{�6w�ˤ��Z��|�l��`	��EL{ہ�`~�^��E&O�g"���0-��X=�>�m�8O�xGB��[�+����9���|���{�U�X�n����2	z�`Q���f���Ko�uC��s�5V�4�n��{�U$�C �k�$G�DRA�H�B�Rq~�E��i1	��z->�����1�e�p$u�<Q 7m�fN�P��xiYF��R�{�R�I�~"=�٪��t6��m^9��39��!�k+�:�H'�M��������nx�lJ�X_�g�g����M�Ek�w>؏Ѷg���ߍ�TYD_l���ܷ&��O���k����<�D0元��d=/s�dZ���Z��A@��ybߣ ���K�0R���^�������3�Z�pS�����[�+_��9�lg�Hѥe�`���*��4���t\zIh��5���%2�#'�C�\�V���M^�O�,�J&�5��$��]��2��w������������ZP�rM� ~v��ȉ�9i<1k Ț��$lzԘ��GBr�������1GJ�p9���]W�8޳m�k����^�§��2�ֿ��)�f��"صe0���3U˰]�3�� �������� Ĵhg�/�bج�G|s�C`�425��e!�Rs��7��
t�'����P��L���?Cp���\4ٖ_��M2x�'��ZY���Y5Eb �j�
g��	S�>濉�f��T��=^.=���:2�8���v"��R�KA�2��r��G�,~oD6Xw����x�0�ty�.�T��G�����=>�J�tY�����][\��lC���UH*���ܩS�� ���Yuv�T�c�=��6��:�����u�Z��X0��V��7M�̉�i�2�F�
f��jפT+�/5��t� j�u���^|`g�t�����/.�4�4ց5��`ٔ�,SP�����*����y�>�L�����	S]�ްH���S�B��h�}b�;i���v͐撼���de��h�R�c��J���@���6qe1�=�[����ػ�4��������<�P)(vl�6P��`T?��d�����3OS��S'��m�L��2�bo�$���lk:�xMh�������+n�,L�s�Fe�O�Z�}Y$���U�L����@�a�	�8�o�1�A��9
B;�͞�#�P�#�Rj�|zG8�$��\��縁��wma��X�`(du`�{)>=�K��r��M�[Km]�y�7^XD&Z���1	j�,|����Eʟdg��:("�;"��%9�'�dn_Y0���4��Ӿ�d��'�*�ͼy��8n�t���tq���7���UJ� �Kv5���:Dr�E� =P뿊D٘V��x�q)�XB�nϐ �\�#BV�g�}��W���Ҹ���P�-7&������W-X��!�PLٿ�e�T٧C��i��fy`66v��e����>�
	?�;����i!5�2T������Ud|Ө�X7;�����+�^���n�uM��M�y:~G�k�3��UY��n�`�����Azݺ4���h��!MZ�h��,n�ؼ�Ǧ����=�#��
<��?_�Ґ8���O�M�^l_��o����{�w�ݴ}���5QaN��1��C��'���5x�F`K��ƚi<��&��PWL
�	mj�V�u�]�3�����fUę\'t��klo�v�
��������M^(������	t��3�>[U�c�z�n�G�,�&��*dl�Q�#�P~Y�!bmq�[<�Y^{fhfX%;���#�1U�tɡ�Z����6K��zw�܊y��Sn[�QPR�_?B��P�D���5�wBSL�Ѧn'<�z#����~LI1S�fՍ���]�;3����3N'W���e�q��ԑ@L��
ye)~,�x�8"�i�|�&'R�#�I`v�����_�T�Cq�"%���D(+�l}���ÉPWA�uc{5�`6�ݽ`��2�qՊ��k._��5��*�*�<����E)H��׵%�j�;�򖙆�;��K������A�.o7����К����9�����U�'��7�Q2���Ғ�]|l�EV�}�@uTy}G��8��:t��h��mX,=��j���g%��P��섻t�|r�zax�����,3�V
�}��N,8��թ ��)�`����i���4� $m�	7�k�*���}�B�� �؋�C~��\ye��ꥼ)K^��)r+����gf֑B���zaWn~�o����p�Y���"j,X6����^��5�Yʽ���~�+��f����~�7-dpg�6\.��e�c?���Uv�@q���� �^�KWspu�f�m��]�;�-���7kؾ�k
�`_>p��+ w���r�o�td ����KL=�,;� '�og��&�@$eE�6+a"�8�r {��M�Ei���"�i���k&v�s%����'�";�~Jy����+��W��ƕp@�%Z�� 7"�����2A�6�.�):}Ձh�;R�&�A~U	� �f��T��9�*/q����)6�)4+��ӐuH�׸$:��������� 0F��_v�Ĩ����=yq
���s�~��f��Lw?C(ʮ�Ȼ���F���?���7Pkp�w|�a�x��|P���%0]~ g��2�R�5�(���̪v�$Dz�<������(0ٽnG"<N��s��4��_}�٥/kd���TS�����&�����Lג��e���$�%�-��'�������K^Ne���l�br�Vy=&/o�G��K;�1z�IFif���&�ș�΁�.98�TpB|eO�>���[�X���j�w�v-w	.�nX��V�v:klQ5Ü�R�W'�k������_TEq�\�L��:y�$��u�)oZ�<���b9[��5{θjڡ�{돭����0a�����g�l�n����v��U�~���~��L0hSh{i�Ou���	���(,7t�@�֋��SO�FuEw8Y��PQ������g�-7�660�,ْ*������i��Τ��ӂ&�~���̺92�>a�t6簤��,`��H&��ji}�0�`CI��oL�� �D��VxX@mK2s1��|��<3 ��{�,6n.���y��]8eI��e�?�>uuA�2	?"��Ek���>��X1�B:%����|��y�p�C�M1��:�a�
?�Ҩ���^}z���>Y��7���6��H8
��Pp��@�)
��������T8����W�Ʋo�����Q�C�K�a�S�2J��Qc6�zViYPr���$P&Ӂ]���56������q�K}z6�wN��bF餘�����o{��.�pm�{L�1':Dl�nԼ��3�"á���3�P���WU�8y\�hx*1z��� �H���Dd�����ڢ�Ϻ�@2��hG�eO�a������GY�Y]�� ޜ����1P�=���̏'�hT�˶taǑ?qİ�W�Ia6UPݦd.١�k�3�<�7�e���B��%X��i�8��g�u�����&_�$�i^ė1���r�R��;_��-���ʊhS�8���	���@����c�E���U{!��lbx�[y[mцTG����~��r�I>��|2�mӇ}�'niI���[rNލ�?��\������ |�=?� ڻ�<+����*{Ӎ��_׈-��o�d^�A�ܬ�3D	=��Ê�F8�jt��s�]2���4��+�t�z�����x�IE���P�m ��Ciw�2w��B��X��c�A��7�_�V/�9���<ƅ���:��O䤏SF/ƿ���o~7��Ò���Ӏ������F(�ُ��@ �t���n�.L�p�*fe�F����{,ʝr'��՘�n{���'��B$%J��Dꮚ (��:����Ȣ���O���-���ǭ�R��A�s=�I}�ܣ7<��-QF5�|*�$�Z�6�=|�M�k��DK�i�_=��(����Ӹp�y$��tr�|�$^��D�7ELS�3xF����_����0��p_��Bo�{�i#�������R>�7�a�6�}H� �V�	
DDݯ�t���wE����z0@�Q���P��Q_���g][���E�E��8G����*ɗdـt�En�Bt�?0T���ntU������6XQ/�o���n�����nz+m�m����{��ȋ��P�Xno�0���s�n=���0�s���3g{�@Jf2�e�6rx�` ���B���Y�Ŭ�1��ٷd,�h�*C��$e�y�Oi����O*;��T��
���+���Bf�4<k�B'���h��o����.n����{�q`���'�\C�� 