��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:'�E�V�}\~�A����Y��?q��|����}PI��hK��Ǆɰ1!��Ty
.�,O8��)��6�N�U2i��˒�]�R�f��G�c����S�S�sv��.ׇ��ܽ�N!��Iy�)���	��cN���@Ge\/�D��Q�K�6������OS�/���r�4��y��f�m#CN5��(l�6͢�ve#f��~��|��U�K;�#�z��$�@����0VT�g)��FRG�������(s����c�}�=ang>8mؑ�ˣ�L&�Ϗ�A���Z�[����%}6��ɫZ�)]��FVhA&�w�	� �+�? lu����$�xwto77��;��"{�Բ!@�v�b"D��{g��5�z���V�%V��P����^e����(�� Gs�^xkXɚ�e�mFد��C��Bt����n]`@����vb��pe������QV>����S{X-��u��P�D��8U1���}�l�A*M�|&�������G��  ZMe0/ճ���1Cj��H����:�Mخ��<�_eI�b��]��[�f=�]����0S5+o���ںZ��(�g��Ǻ?&���=lX>u��6n�.q�V6��Ga(���̚�A�[�pI��v�}��;K�w�B���#ڼʌ-g��r��$�y�����}"N�v�H�\uL�G(,n�����ߵN�r�ω��BU6�����V:f1c!�>�̻��,�1iED�(���ot�f0�\����TvWD�s�	2�ˌ����և��5��FC���Z\԰9��@��fi��i^��.="9��j]?����l_�I�`<~�uj�
Ƴ\v�l�j�������� �w�3 ����t�.66�j�:�Z���*�Va~�Z�v?��8M���MD�����n�'�|UN��]�ίߌt$��C� �)k2���m���	o�U��`��T$:�h�.�	�����;��'p|!ƓU�-�9nA&ԯ�G�n'�g]��=
���9�P���	8l��=AFeƍ�0J,C�n��D��mU��<n�
�9ş�	Co�y���!aʝS�{K㫠06V��{\$��l
�+"WB���v�k�~J؃H�^T����R}O�r��@�N��,�oG꣫\f���@� h2�K�3b�
J\~��i/����US�¶��1%NS�h23��9��|�y���k
a��.��$���d��=dY�T��.&��a9.�2���shA;
��e���8�����^�ޥ�
������9���`�����r�L�H�\gCHCe���Q*��7�6C��JnB��ɴ��lXW�{�U;�k����d�"�R�d���ݸ� R�����p�
��a�ZNQ��zm�-C��hbc�F��^b��S�C���PҌ�KmL��"���F,���J��N Ձ�4)q�M@���堓k��(2�^�4m�
L����u�uG��69Z��r���rY��YxX�cZ�#���"���S0|#��T�����t��;���X���� �[��o�fS��2��p�����B���")�c�7�r�	+7�湯�q�MY��To������;Յʇ���)^���0#n����A�ͤ�𮰬�D���<��Bq�K�Tȼ���_O}���K�h�=�g(ZF����$ރ�tl�Y���u�u�V�i����A�m�����U��c�<8�B��a�p+�a\)1�G6��&�TC��T�o �Q%�eV�Uw���h�8u ��2�cWՖ��y�.�8!~�#7����]a�� ���B[�6����ʸ��u8g/��`�ڌ�)m��d�A�I� a8�Q��9��`����t�@ZzԚ�)�LCw�5�4�F�н.qP��g܌V��$OeQ�|�ȶv�<_��a	g+`�� ݿ����E*�1�U�ݖ�|���DS,���}M`�����.�|��301#4v�y2N��\ׄ-?br�ÒX���.�ߘ��܉�;���:�S��1ԣ�Y�X��5��=SťC����Hj9�����O��5��0�l�]�������D�{��\h�(�"jK�}�������IP�v3��r��\,՛ � Z����h�Z�x�@�hK;�޲�A�:��f��o6@dWJ��)B~E�R��|���4*�fQ�ƕ��X��k7�(:=�r����.�(�Q�˰ [�ɇr��#��%���Q��¨L�7Yi������d��(ŕr'���z��L�8�xd�7�7��s'��c<�n����`3���8�@��������637컅2Q'�=�Ng�����U8|K9zX�����^m�xsf���S�	�:��St�a�D4e]up���< ����L0!љ�{iI���C��B\E���� �\�A�fA�W��k���a4ChOC�'�Ξ�� W8�M#�b�7
��x]׼ $E�A4���&/*h�{	Oi��򡧉���[�����,�scD���!"Z�47��l���k���o~�5���v��7`/����E뭡�����A.�|s� �7K�Az�c��p��O��u���Pl����M�z��!�>97��N���Z�C��\V���PLю���� �Lk����|n�
���R��U���]v͏@��wiP�����Ҫ���>�	\]�Q�4�"�Y I�#�\�1�؏bˬUʻ;FO��� ȿ�WF�Q���ՇQ�f�s��P!sjI&�1^����q �N�:�BpJN��g��)�$�a�EIV��y�	�O�ɏ���Q�/���W��?ijT��f��K��^)K�� �V�׫��Ѫ�!�ʢ��TRp�Xtԣ1��d�R�����&z�!��+���%��;Z�À(��H�x7���n"�`�� �n��k��^<g�����u�Ђ`Q7�0p����ڪ;ѹ|Ҋz���	��/�.�l��B�|F{��IML�J��]��$K��4ޯ��	�A$�Ս.@.� �]�a�kV]��f��'O|�a�H��q�un��d�\&?��*�R�?7|,��ι�:�|t+J�,�Q�&d�@�M��ޞ O�ᵱ߈b�Z�l��c�h�w��/ȣ���q�������R�+�w���=���|�IEA*0�5�X��5�̑eᯁ���'�";4ٗ)�%�qE�~��nWV:oR�ْ:)���c��y�q `t�
�>2%c�Qt�Q�.�l";w�7is<�-�ɂ��?��Z�*��K�4��Y���d�*�/�!28�����&���CpO�Y��L� ؒ��u�'������D��b6�!|n�����-
�C�+$뉐�<�����.�����vb06ٖ�TTQ�᫭ �7dW��d�d`>�}6�O/>7u��	�ƪ�`��2j3iT�>�K艞(T��p�}�U��ފ��F��qs��|-�ƸK$��f#x: �5v�*HY ]@Ԕ8~�*i�6�q�Gߣ�hU�@��8rOB.nW�TPIǐ9X��&��?�Խ���v2����.��"�j����u�
��p�ς��^`P�G-N��&_PlSD � ���n���8���SX��2�}�W;]&��Ot��)u���&�1����}�����(EfЗ�*c�k�d|��r�oi�1_��[C�d�UibI�yp�5W
�F.�睨� �n2[�4�k�c)ɍ']TW�P���3#\����&H �o$ї�F�0���~ZY�I����o B�� A�G�c�D��SG�|�����'\әն���@�4�Şb�I��D�mb1�lzo3\�j�v�Bvo�/����m%{��a
��ѳ<����;e���LZoħ����u%F���=BƖ�N�bkj���0���[��ILQeɬ�%�(Hu�7�Jˁ�j��b��&9�\*I��|��)p	T�J����J�[*|m2��h;y)��tDҽ���'����S�)���S�p��ײ��⠗Rz�|en��7�J�Y�V����3-�"� ��wv���jp!!��OOgV�X��GY��ҕ(d�0��u+���{�~+�&��|E���.q���xPv�7h���Dʐi�h��b�`�]6��̕��>���MW���6=J�3M1?Č���'�t	YI��[��
�)�e㝌k�Yz> CC�`Ij6E��"g���cv�]!2i�W�����`Y|�yC��AO c�N�]�h�\��6�ge+�l�;H(����^sU&_�Q�?�1��:����j�F�q�'�j��+�|��4�;���G���B���u��3�܈ݻfD6C�eBb{`���y=�"@��~�g�)�������O�
R_�D� y���`�׏�g DTÂ����ú��ŀ�V������e�|@Z�*gi��⸖����l!&������e&
7D���%e��b����f!�x��� ��;D����o�����%[����ܧ;�8�`bh��"_ey7���5<��~#+p8�k��-T״}��Sr�	�c���|�f�ُ����;>�%��5�KsWM3��<c�_'	!�M����O|p�NS�χ���=�C�Ә"	Y�NM��m#�.V��0
�ݔ
,����0̬-#��%N�s2Ǻp4�P�$LՍ�l(�}��/X���ˎ;=�)��K�Ȥc�w��k��v���y!�����Vd�B�R)��=�����
� ��� x�Fx���eU�_��s5S�Φq&����M��"W�e�25g��˻gQ�"�\U�+���l�MO������E#��st��C�躞nc�.�OaH������m���(Hh��y�q�SU��%X|L�m��0K�VQl�$U)���7`2��0G����d�Ǐ�����g!NU>#�t忟��4� ����aH`�ø
��QQ�� �=q����]���a�y����3�F�ز��Eq����t^�����@����Q��=@���pԾX{5�� ��n��9^>�����Pm��:�f�P]�A��LV��`$X	K�/�� ����c�S֝`�Nx��^���D��	�L�ʜ��T��]���2�
���JP���0HV0x��閥/"W�����mdK�W<w�>>+�[W�8�����ˎi�H���� L"���3v�j�׎���Q�~�����T��=�8���_� ��)I��a�%jz�;̷�����6�O�'��tS��q{�ѣ��cCy���"��H��ls������u�R�C������!���y%�Vx���!�iJ��6 ��{[U5^>�sZb��T����pФ���BP�,��!K� ����7)䊤Ryį�Ē}�
���7�1Qe�k�Z��ogftz	6��`�U���Z�GO�}�~4kT��FAL�k��p,J�q��[��~$�S��N�\A��&�;X�	��!�R0W�9��זU�q'��~-Ҍ�ၩ���]ƽR��#�g5�/�F�O�U��6�1�y�wx�z���g�xi�r8E�u�ĤAyҘs�O�keb�[[+8�>�|�s!O���%�mE��[��~��˳�Ar�C�����hPO�}� �)��1����EN%���ڀ2���z����w����Lטk���?�>/]D���-��a�24���9H۴�'Oc�����v��J-��5B#�23�����8��Q���Z�j�ݗf�+���OE��q �岔���"@��v2�=�ݓ	_�f./�����jb-��c�yzM��j�&�������8�(�p�T�Ӫ���F����j��4گ�Ks����~��aј '�-��v�/;��D�V�e�a������c��
gV5Dc�,�8�O�S ��(f�mR�`S����RU]d>A�*� �Os���ģ-���#]�|�җ�ڱ7��
_���%�Q�_S�����=��Kx���Y�_���%p���d��(/�'��t"	T��9utU~=q����c\ws8�2'���y����v��s���!я�og�H���$���q`�S�v->�@���A�v� �d60`	$3ijl
��L$a���'���`4xmw���hZX̾
4�n�a(|�i䬪�cL�6X�Du�s��.�h��e�E3���:+���G��ŷ��/�����-8+���߅E���'����z���1mz�I>��N}���FmE��h�e#�u
j&9�k��E` !zxg������,�,A����F���fJ�n�:4R~��4�HlHp�'bT�i�RA���Wr%�=� 1�1�@L���1zD>���~�؄V@�%<�MY�D#�G8��g=�"8�V�p�'�2�Q�,o�����6�KL�K�;��]�	�g*��i
��>����Tbq� )xٍ��z'p�-�'��,W��H'�=W��U4�3�\��X�ΐ��jc
F9}�0i5��ƕ ;����	�pm���=�C1��a:I����p�{�;����{�o'�h_�SJ"�+k`����<�3���7�˩v��E��ۛ��T������t��!ۮ�#t����!H�h�M
&2a��R�A�q��ujn�Ŧ���Wu�WpKi���j��y�Mgj���e�����ր�w�d��G��+���/-���r��gl�%n�G<�Įl����#���^&��|�f�s���&%D_��(W���M��=b��sF�۲}s��z���^i���(�봳��8	��T����MDp�^k��q����=3i�.���-=�#����~!�2�J���"�21�)K��]�T*�B�q�#E�k�R0��P��:��G%lv��������(փ-�K�JH��<�͓쯠��a�L�%�2��F,�T�'�r��Wk���q�UD���r\YG
¶~��� �����K��z���%�e���\����Bܹ9�L<�r��Hݖ��QT�_�<Ҿ�i��4Y�� >Ws\.�$q�>�Fc��SY0�訊�$R�{�_
\]�9�1��y�5�P����v��'Hjڞ���5-��khr��W=�bz�-��*��v�;���!�D�YY֦��/E�{f������b�"P �%urʊi0���-��S��}n�6�;Ccus�yŝ��s��dj\���)�?�]��t�1����� ZV
!����`և����)f1�VTW�S-%����u|�1*�]���'�L����S���܆��^�V�R6(��Cjm�H^�Oوv�f�/�V��%�|S�y\��S�a� ���;�&��5��~�T���X�ZY4P���z�P���9Ljw�|��f���$Ծʁ
��d�*�Y�?R�����XD�=��H�pT�l�k���sU��B)m(l[��߃!�S�aD�]AOX�5RU�Ѵ�*7m������A�1��xE�����tV=ud����f�y�����{�x�� ���z���񉳇rG�G�c!�첨Wi��п�H@�]�8�B�n�T��Ө*s��K���gꉎ��	>�o���
A�����N��r��ߗ�σ��,�4���.�L�N#U,���yJ�6�Ox�,wB$_�j3N�.��1�]�d�r�������I�ǽ����=@kUnLc� �%��F����sң���X��X�8���	�Hz6^��p��`j	Bόk��"��l���.���?��&0qgԿ@�t3X'"ܮ�� ���N�3���@f'���1V���(8��.�e�@q�uOJ���_A�,1�$��H������?3D������F >�Q�_�(�]9�� ��N�c�:	�2���mĔ����o���ptPyZ�Ҧa�D�#1c0d;,Y�Z���$?N���vr,���A9��!(��R��ہ���D�c�e��.joTf�/�բ��jxo�,̤��j�mMd�t>}�O<��O���]��=%�	݋�s����b, �
�%�s�Y�Rs0������zsgi%"����b=�!�����o���A3�z�=�C�b��S�v���S���Z�n'����:X�mm����
�\���3�t F�mA�&}�>�kJ)�X�����������G_5,�>޶�N2`��=PC�F#�%�[#4��3��B2V�~6�g"E3D�F��?��[�Mq�C��u~�&�[Z�gy�q6���2>E�ԢB��.�/i�"�WP&HM�}��j�w�o.煭.�Y��Lp��<�疻j��m�b8)���S ���S����H��鴸�S�B�*��-��c�T�A%��)��\_ ��߱xa?4�v���6gG��A�f��9���I�h��K�����s�JqfR����)��5cݔd:��5{πܭ�1vf~]�ڭ�-��H��*�"�HJ˴3����ȗ�h��8������OD�Km%�T~H�îU����b+:;��d Kc������zD��?ţ��y e��*�� ,��{��8S�i�dC��\Bq
��x��M.��;~~�������xݻ�zD�#�U���ά��z"ę!R�'75�V9��N�49?nǽ�1��Q��R؂x�9l���P�X�Q���*�UW��X�RӪ������ՍC��M_!�i�$�2��%����� ���1�Z�Ud�˘�!w��	�\9�2���n�2s���#3��Z�-�Ӓ0�q}_��-���{׼m}s�7ϖw�����IN�j��u��,��P�*�����?�a�q�bv�I4��� ��n�&IZ][L��*��!@HјL����"enp�|��t��tX���I�"����@�,uv�k�6a���]�A]Cm1�������bj�%yd�0��?g��c?���
L@V�<������i�e��4�t.��u6���3��|���Z-e ���'�n���q��)2�xna�,�lR��(��z��A���l�e�/�ܟڪ��IQ� ��$�V�2*�T���v��Ε����8q��*R�',n�vE���|��ے� �$�a�]D�������&k���d����w�k-\iRi�&�U}��=��ċf:,!��5W���~�j"�wc��t�7Â�F��:��K�}#]��2��N�
"����ᠸۜ���6��W�&�Tۧ|�.�P�l
X1&uR���CbY��䉟�=V+���sZ���څ� ��!m�������KV�q"��ҵ��A�$�����ΡW����yp��k��157a�[��=�*o?ٲI�U��$B�x���"�-�>�Am���vWy!q�(7h3Ks�
k�d�4N�WH ��k�A.��jZ�u���e�s�*l5�G�4|4�rWK�"�v��pQ��␹������f/ ��M֟��MW�+&��HQ��zB$�{����F�g���x��Yr�M�J\�o�x�c2k��%��G��yB��s���iA|�|�s�P�~W�M;�=͏w���P�Ĵ\�HЏ>Y�����Y^:#˞�Z�I`�=�#@O�9
��&X(�*-�	;4�҅�J.�E����-l���-��
>R��]*�����q�,=�-<�"��%�[FE��(c/�n}!z}�i�h���8���V���?R.��EK��<�����%���H�dV8rU�L�b5��{�����SM����M��X3�q�4�Wo{'���G��Js;oq�[@�(�8��*v��_U�iB���>fM��D�u�[���^XK����S�X�9j�!�I@�I͝�gO����1�g��R�K�:P�3G�Z����P���@Q�*�y����O����M����̷]oJ9���R��WUr�K	Э��U��2�'.�>[\M��������Y�ֲYx�������!� Zqfi�˕���ce�ǖ�	W7R���p^`9(�
�`:��c.�I	:q�%ڼ�|�+�Ip� ��׋!���s<Yb`��oX����QȒ��/
}桠���V��ͭj���<n�!�5P�ߣt��>t��ϵX��۪�*-ڂ@o�,���t8�i�r��#��i3��);[��v��-]�0��L��gF�A���+kvs��JW��-��ho�N2��D�}�ޘ쫟���qf-QY��>���3��D8bh����EB;z��rS�d����ٜv>�9Ŏ����+��0̳�n[�{Z�>�H���݇�W�3x�EP��j�M�䔪dM_Y1���,4)���g�>=�#�L,����"�X�I�H J��!c�_7�M�
<�7��/�/�$Ή�@@.�:���K�cࡖ�v^�Y*���\�����go��e���d�����Ry5'p��tk�}�	{W��MK9�*��U�GF��#C���^B���s�C��vUW3l������$*��z��IZ�y���-�R�T� �v93��v~�NFＺ��Z����e6WK����D�{	�OH4˽L��������-��9�.�>�:ۮ����d߀�$�����\a-?%O��#��>�c���a���x��,�m��/�Es�2�H��IA@5�L�
�>V-��ӗj9"��.�sr.}g,��<�ӪnU��'��8ΐh�Jp�a7p�����i\tMk�����k�'��/�6�${� 0!7���2&�$���i�OÚ%�%m��S��]������Cl�?���n���?,�ej�Y�L��nI�	�B�n5p6��3�tv5�u�"lj�7��ui˖s��W�4**�H�@=�&�Z�~����c��Hb�������9�y��$+#�=�O�8ӌ�#'t W�L�/b�̑4|�镼�Y)��1��i#n��(�
>�8j�ԽXi\Ok�%�ؠ�(s�6U � �K�Ͷl����{��Ћ.\>Gי���e�r��&pr~�����i��*�*ɻ�`�%[T�Q���A�+EUe���rz�.��ՉM1,CS�TowHӗ����C�mQ��̐K����e�����f����OU�=������,��=���4�S��t�1 y��?��c�{<r�ծQN�}�q�mZ�UӺ�36$>?�ҕ8� �q//���>�$�|&j�Ǟ)�xXUu)}�o������W��U�T�s� s�Lr 3m��N� ����T>������&�����A	ᩊ3.�?���D�\o�ݜ?�b�˗���W��5w�^���$�}��F52E�]�S�V��Y���H�moRb[O�����A�!��6�[|�b1��o��L%�0xa	(c���"��[���-���'�{��7���L�0�@�x�?/���]'��־�[���+d�؃66��^6�w����cv�)�2-����T�\�/�{��e��0e"�Tz+�Bݘ;�ն3��|#�>`�㞉�}>+�vV���f�&�_L߻o!�S������� [$.#��4���+�K�ي_9�1G"�1�9��5ff������ǡ�t1�k<���8]ؾkQh�W��$E�{)j˓�'�br�M�x�*e���p/V݈0���<A5^��2�w<V�Pwƒ[�I�q��ou)3��j�{�w�3+����|� �����#�82;�] D �N{��7Sn�9��XF�W=��ꏰg͹5�s�IعxAN2h �Њ�:��6 �)��ұ�(�w��C�� ��6�W͎�:cԉ�����~~�r��~�F󹇃����l�$�0G��	���Wgֳ(7��?oP�{|Z)S4-Y����2CҠ��I��!
�H�6ؐ9L4�o.��sZw �1�}������JN8�mW��,��qu{�6w�2d0U)��XH�A^��~a����_Veav:��V�T�q:s������H���ȧ!��U,�f�T���i�d\�]���Xւ�*FSµ�i��S*G{��j��N��!r$ejY�-~b�3W�8�ַΉ�q�lv�0��4f���������HDT�!�}D�Y\�k���p�@�T�I#Z&I�&�<3��-4�����L��<��G��1�z�*�eʆ�a��.C����c �@Eb̚�AU@f@��	cA�c����ڙ�B́P�N�D:��=�6s[.���e����;��gO�p�r�vb�Ǉ8<�l?�-�f�<D��wJ�q�[�١�Y��Ȋ�*��A[B�!��y���Y��n�|0�x#-g���Q��t{��&3t`������� ����Y|d囫K<����K��p(��N˃߹-\w;尻���V�s3�	���L�,&�p�_�Fj��>CX�h���R#�n�ܮMՓF= ��>��h�MqwU�&��� Eʕ`2Gjg?C"d���U��|�P�}��̧0������]@�Ùܫ����r���p�������ׄs���?W<܍6R������^��4qe �L���Y!̝�h����7G�W��ܥls
<+>ȴ�`�K}��њ?l1k;>�H%�_;����+�wa��!ZJtJ�s�"h��Qj��,pxݫ��m�b���O��/�ǁ�]4�O[8';\��%���kwl�xW�i��rymǫZ2�Z�2�6!T5���ҩr��H�(�kd1ӏz[OVV</YW�:���MXjc��p.G����QO#�m�?L�ú���L�e0�H�چ@��c���r\�V�L�!P�ھ?�/1ZpY���B�R��|y*���
����-|j	߫>3�ʍ�����,V��M���߁����I��y��� p�y��5FK�9zpv�����C#
�̮m=!-	^��OP�>���� ��=t\��W�	@AG�@���5��c�[��.��뫐*~����*ҟw��O"�� ��O.k�0e�AƔ|�	�H��uD�$�ؖܖٔ������r�#�����@[��sL�����ŻQ�g#2*�ѫh�P, }�"�vSH�)�o��g���&X)a�V�U�r�s`�b�R\rk����Z6����S1d�I�[#���T��?~/I������u�Y�G�T�Cg�S�����[�.=�{�0	z�)���ĝ��K26�^7Gk^Ң��h�A��E�6�.8���.>����蟦@�i�J$]	d�b�1]I�*��S��F9�1
X�.n�"��yxZ����IU�ҫtr�qïu��>��2�� �S�e|9D^<��Ote[�!wnԿ}ZƢ[����XE
����yۘ��#m�s�׎�@r\D�K'+E�%#*�3x�%1>�<���UkԳ]�Ϫ��&�Ш�8�Cd&������p��!#\6�{w&���b:���|��2��Kϸ�Pix�MU��nĎ������Lȣ���Kj�LӖ�Z����_���C��3�Ð�Tԣ���Z.8��FF�aZh�D��m�h�+̉#���?	u���<qD������d�qJ8i��pK%�����#��Rve��{�C�����F�g�	������V�X*7��#Nͤ�JeA�����6�;�E�����@�S�1(Uv�i+���ub=�Qٞ��K��%���~|����G5��Me��,�[�J��H�Ѝ�&�`<���Q���%�B��t{�GA�ę:
=o�:1ap�1�l�s҅��d�t��3