��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���yE�42i�0 5��l�R����꨹<ڛ�\ �*�L���T���DL��3S&�dC{��$�d���T-(8�n�2����L�*��1�8�PJ&P:D:c���*(�w�]���4�x���J-�h�ҁ�`�щz� ŉ��Õ8n<�1$կ�����鰱� 3Z=�e�7�cK��K��F�DE{�!�v�:�":l��:�b;?%�}�5���p��yH�,��*�h<��p�)Q�C��>��=�?����} q���T�Q=Q2^��0Q��P��'��t�R<�k7�6��F±|�Jb-j��Ǻی��r���}��
�)���Y�`_�A�kY�{��>/Y6�
��u�4A�j���ĲN�ޘk�V	W����ݫ��[W��
!0���b��p-X����aF+DL��+��R�(#:ڋ�����Z���v"�9�������BK�f�d�l�2A΅�z��-搾��,��O���NqK#+j�W$=r�J�ݎ��c���25q(�Ld�$^�F5�O5]nc���e6u���6ի݉��˛�����'/���y��a�nB��	Z_��t\�X�� 3Vu�G�s�7w�{/�)�"���]�<����([#�x�/��>�%vr-P]��p*�6 .:'ɕ�D�o�Z����&�P�b�,~�v��f}Oũ1��T�2x�4��:���t[��[UP�؉����ʓs�M�S�K+�Z5��`�+�Mm�I����D�G��C{/ɀh{OWߜx��V�v$�G뛼fJM�V���1�}:�Q�z�n2�H�U��θ�{�6Tp;p�ؠ��+塖$ol��R'>�hm3�A��G�zSmf���#��:�0�$w�98@	��?n	�l�D�Q�I.�'����ÊGc��s?���/�ۜi����-Aφ�jc '�t.�L�(��Ȱ�a|�D����� �&a����D��fbVrB8C���`��))�"��VC����&jO�������i	���%>�@��#0�Ӂ�$՞�$w��0��Q@�$�G���i�z��u
�r�}]]�\ˎ���E�����$���F�+�a�Q����<%A�͘���~���ݤ��ˊ^�~E�j�ʗM�u̘o��aO��ۓu�=G[1;r�eC��>&��b	� �J���-S��=*3sz�R��$�}��X������Hܥ m�k��hC�L��=/ٽ]X�P.c�G��?.���T��X̦�?	��Gn4�ЫzG��ᩝ9O�lxaW�{�βm}��
�g��d�9Y�{�6��ae��Y
�a����]��f�ޚt��f��.gH�tN]�	a�2w���0� TF$H��x}�t��k�_�&#[��ZrѦ%Мi��ׂ�k��f����4y'���;dQ�䣏�uFv��o�d���HQ��������~�J�t[K4��:WJE���)8���zF��jK�[����$��f�-Dn{"Q��Q���c�������u?Nh|�\��/V�����Q��rӬ����5����eSS�	�Ԃ0wͪ]/m�����=�O:I��?y;J������e�w�"տ�M���h�؍��k��5�o�J��Ľ�l��M���zHfq�0�0xO�@Tx�q�������m�e�n���o�$v�EAI�vWF��/�t��W�MTѥ̄��z�KH=�
M-D���)�B�ʹ��:��W
���K�1���C��2���3
��VRE�"�D�,�XrAB^qRI�V�E�[d��,�����[��m��$��>�]�-v��:�Y�>N>�:<��y��ѭz�,��r�"_�Kp�1�����a�/?�v8�𞿀3G����7n6���Wظa�������C4�.ޱ;( ��{%����� |N��Ĺ���gG�U�2fP^���CfMJ��T�����kx�Pc.+��%�crm�!��n�$vd���zY7U��.w���c-����<����ߺN�Z��Q+c�\���B�61����Z��Qܳ�@�>�\��;�����dQ���{�M��;���}�9L����F��R���0t/�V�-��(E�dO	|�4���!���p̪U�`պ�"2����*|���N����MtOi/�j��%HY�����G���3�S '��o����u'��ߍ��ͩ'�'a�iO��	�����_��wTU��Z5´뎛(ܧ��(���'�s����_/��� BB�?�;<�6�J0>�Ѩt�dQS��T��=�ua�kVFo�l[��
J鱴��m�:��!�j��m^�n�.�\@�m����l�lMoEgG�>���.���4"�[�M�v�Ѐ8�O;ܛdI3���3��n������O���
�z1dc����Z�����+���V��K���Y�l���ޓ��5�\:yW�s0z���Ms?cW*X�M	%���\�~S��\vڝr��i����FPH�C�v�bD���т�K5�=� �j�3����}���7�<@���e�����H#;��l�,)Q�Q�r�+��^�l\ڟ��Ao���������W�l{hy�cz���0�h�V,/�yhx��t��%9�\G[�j�ϑ�e���Wy��	��W�^��o�t�p��XO���
>`�|�FP  n�=[4~�*���ZsD?=wF�_1���"��i�kMpJ�$d���L	��ڡ��H4��R��O�Q���yu�{E�ə6�CW�j��:���Rm�*|yCȣKsQ�ˇ.	�~�v�R��ںJ�t�qd�h�9)��	�3і��j	]��/9ô�@7
�*x'C:��jBj	�+fYY�px"��6�cQ�0�M�:4���"�5�@�T1�����U_d�؝�65�Ω����M��:Dm�1���6?"��|+�#���:. ��᣼�jDv�װcе���)R��k�_��6�\~-n*T!��M0�G�j��Uꀚ�%�c��� j��k��Bw�?�ລ��R�P�.C��`�%4�ZQ4j��.r�N���O�I��ؖ��sa�3?9�YFV� ��![/dg{ҥ��%ռ�o���g�,֏�!�P�'d�X�zj=1rL�~֬�K�%����GY����!p�z�H��S���;o���1���
-��|��36s���侅d� G|yT��Fj��N+�i�b���V�\�Vӿ�A~�r�w��nq�������{���-0_�N,�� ����;7�'�'1`���D����^'�,����j�5��%� �����@��Hco�x���|��@���/ /���՝\�D�C3��Iv��U�O�/"�	����*�uW*'�3㔂�gv�YN�L���Ւ+Ƭ#�i-J6�,C
�ؔ�^ڱzN��x��}�L�l�	���*K��»�AB)t�ڄ#� ���[�/�M��N퀹]#���%����O��"���c0I���p��a��J߂����2�nΡ﯐<�ñ�W���u��c��O~mP��	ɰ���d9�F�#Em��,��)��m�
 f���ʈ(U��DL=�ˠf����`�H�l��K���jڱ�[��2�������.��L3��2pmǨ��]h�����U�1��-9-͈[3(��S��Am��b��H��;���G������n�oiFT��YT2 ��jN���(E�.�	l"��ѿR��.�0~��w���̲��(B�>R�X�טb�����n�T�����H�qd@q,�՗*U�HuH�.gB�.vdn����YF)Y���S��|+l($;�C��M!�ʙL>\����&e����I��=�*s���y�鲔� �$�y-3DGB���1���F�8��þ|eujW�f)~}CO�����tKm@��>bΓ�`T�Q~���	��k��B<��m�	iS��ɐ��<]	��olZ,W]'�q2N�u�`�p?��8�]�v6������G�&<��E��MK�F���-�L�� �c�Z#��?1p+���#�D�3����77u)��Y��7���#7�k���m{�3�ʇ�j��ڏ��K��ϵ?S����[�Lo��%�D�7Ȥ������pD1�@���_Z>����)��{�k����ocB�˪5+,���%�$BL���NBB�}\c��ά!��𻊇���_���C�	��=��FhnV/4��a��QT��e_�g��0$�T��g+�W����������T1�͢�hȌ�9z��BBq	I������`$S�^�����R�٭�b����CJ��Tct@�u�Ve��Z>�x�{�jw�{�J>.e�?D�vk��ox�r{���)_���E�haw[Ҋɫ+���g2��Z�۳rQM�^�E�)�U!�Y�Ρ�^+�f���a��b�~��0�� �ӁŒ�.�x#Ђ��Md��U��7{�2L������FQg�n�Q�bIy�����3U�}M���m�z�����r=W\��@�d�q�^z�>9=�	D���Bt�wpㄢ&��px��+��]�'��G��Z�l�
�Rj��@q�݅sz�1N�_0ð-�c'B��0)`��k���|��j�;
\��:�����ISw::i&��2�}�r�*ϯB$�]�fG�C�Kv�J��N������lbj��UI2U*��B;?N�: Q����g ���s%�*�^�Q��)�����H���9��a`�����_ڡD�_0'��uf��Yљ���9c�s5<`��{����<f�����6z��ǒH��Fy��B3���$�o��������2S8�3 ��D��F�^����Y��]�Dz@��twy�q�O1/\�4U�ҙ>eΕ�;G�w���`]I $揳�����I�x�M�j'�������ub'�\ϯ�7�+�HT2j��qM�lvP���b�՞0 t��8I@�¤*'} r.��Ck:�x���^���s ���M&�%���O������]�=��߿H�����q5�/�q�X�Cx����2���.ne,�#1$z�E��:iI>�H/]��[)t���X�o$&�o� d9e��b��-h���8)f����Ӄo�����)X���`����[p���ȝMuN��%���q$�f�ە���P}��ݚv���7�2�0_��|[
������f��R��6����K�x�E�+���W�����4���ZZ��iL7/�۪���m����ש���V��V�{����6 sL��F��8�CAUے�{��ou��]��b�rf�=�KI��-{TV�TA�D�'�Q�{���h���삀"!��T�S�����]���yi�E��OS����D9�X��n��aw�'_¢;q,��a�:�K�ȅ?�����G��)��g�����4AE8�Tf��n��x�T�� h��G�ܧ��F�&�9e�4i#�p�l�� �7�_���mm��`F7�C���(^�L �>�2����� ҉�9�`��joL����۴�E�<�4�ptH����H׃3X������
 W�>��7G���3�������"Z���BƢ@ܽV��(�I=92�tv�Ӂ��P�J�o2���wع,�]�]!���$��4���o�Uҙ��C������Z��\&�>�P2b`�V1�R��q&��$�:׽W�ȘN����]�o)M��#'S����#���W�&���xZ�0c���y9?P�������mҵ؎��R�K.��i��#�L#��\�S'���4h�4��l1<�����,�!&�|�OE\#g����]����H��
".�O`��1�b�7on�:�X)U+l���n��[`ש�q��B@���1�\W�Z�l�7���k��w���<����s�~?_��E���Z赂�  "�O#pxaLDi4����'b�W��X#c��,a��>�����J�p�Z�|	76E	/#�Н�9|0�oS�W�`{��MLʌ��e��������;%��̇H(�R"��j���,�[�>78dRA]9�,��N�3�4Ī�F\I�`n9Л�bA	6��CM�uk�5(�ڟ��M���l���`/�;���z6=�!�c�.E"��n�^֟m}��8q�q�_�|�� �$�9!4c�a�`
ƢPư�F�7�?9�6~��5ĵ�s�%������[���j����^1x�'�Ý�R���Qi��&�h�èI�(���-�����i�o�$ ��1�a���%9�:Tm0��,9"�?z���ԋ]��Q(��l���P5|]�0�>��:ޞ��rtpꍿ=����.�ǂq~�^��w�6"�4���� _�I��G���l����&XP�*DK=�ڬ?"X�?��jLd��A�]h6�J��>4U%p-?�m��CS�����њj�xNa�Ɯ<���s�Z��� ��2܀Qy^"�%z�e�+����3��� �.喔,��6�J���}]��q����?�[H���.3�3@n	ڲLX�ک���Q�l8��w�c�������	Χ�C�0�9�!9�5ۊqE���|�2r��������S?R(���At�	�@�JC�K��A�=,1Vu>7�[�O�
�{��ͺ��i��c�������/E�|m*q�J�"��	���T����D���{Dۆ�4)#F~�O��A�8�-��B~����<@���}�-�{���=�����/��	�n�B�x��7~*6�����!u.X��6���v���L���d%���д����_6|+��NG��8|��
艩T��R�ٗ:�b7ˆ��V�D2�>^�Ix���:�k0� ݴ��l%�=@ą#��Y1AP�땜�"��ѯv2���;׫���+U�gYx�6	�]���u�i���v�t�QwZX�/o2Y����v6)���n�WЁ˚����(�l/���V� ���C��ߎ�� ��=�f��d	I�0�n6G����$����B�/޶P�r��(���N��p��GDOCG1�H�������A�����p�2�Z��=>ŗ^������+]a�>S���weM�g�n�����C�6ܦ#p�1���m[6G���ڍ�#Wp(l�C��?\�>.���П�.�	��BP�k�h~��v,$�[x5�%��՗p�M?WGa�A*�-ϡRP8eq�q���~{=�2~0<����*d)�/t��ֲa��fAa��
�66܈���nȊ=��ҳ>�R{t+�HY@�q|��Fc)}�m��G��(����Vk�P��OQ�`��,	 ֊�?M&���4�L�V��`�O������猁zl=<-ʒ��d]�K�Q]ͣ0݊��G!؞�'�Vլ1Qk�^E�-:p�i,��{��q@}B�BC���.��[�DlT���?�Ĥ��_��X�!Oի3��33R���m|����J�:��m3����a7�ÞXq&�ٵ�y�[�W���p��J��K��Xz�kq;��3��Κw4b����#JŜR8v�A�c��}2��g(U��Bo��0(	�Ij��$�fH��i���w�����"�b�%$G-]����^G=�fu*�W�+���)Z�~&�J���ه���7���t��<�4��~�M��J]�yJ��.\w{��
��%��h`���	���-�0o>\��)��v��p��b��:��>kI.ʅ{�r�QONKC������b
.�u�T�T�[إ�/��ns�X�����E%W�u�L�|	�=Ѡiw�$����i��r¨�qXOn������>I�Q.) {�3\:����x���|��&�.���}&^3���r	c�����-dM�]�SU��O=�`�ՏS�ҜH��Iu4����UI��to������& >��+�P��+�1��17b�d1�h�6��[vab�D���A�5�<�}sHs�C$Zf���%:dK�1��2{&��6���t�sNH�<��bmC.�l�2
��|̞G�\>���F���!�]���sL#(]g��=R�{�t���+�3�k�Toh���\<���Þ&�+�1{�1�#�nl+��F�+2D�/<j*Z���U֩,&}�Ď0�KΜ{�,��b��BT��icD�^s~R3>7j��jE�(�5C� ��~]+aϔ�`z���p��1<����ʊQ��ӌ*$�*��^���*����'�WR63��|�����F�/d��"��L�C��"ɤ>�Îk�Z���LIN4��6^`�n��)��:�<�0V�+�X�������3%j�C7qY�-�YӏBF�|����L��g�����S�&�?�F��S-�2Q�=��ω���ki���&Kߛ�9$/�#}�:@ n����)&�����+#!��UĦ.oj�d/���LxM�j���I|n��D�p.H6ƥЏ̙���}u��WC�
#fE"���o���� 	�zŎL�ʣ ��a���R����X�/G����e.@�g�[39��%��� ٠LEڔ����R�﹚��P*��v���~T ��j��NY��+���>��d����V�S�8 ��H=�a��D�A���bJd�^k��ۊEw2��*�ĀTBp�}�ȧ��^M�fQ�9�_t>͛G���?��Y��Lge'�wt�x]���dh�`����g�����$��V'ò/	dYC/��=:]vd��7�/2z>�]bG���!���۾h�4��{vb� E�m.U���"��#^5��	9�7b�BrV�2�NI)z{'{s�P����1���t�jS��*L��S����=�����8��5d�%߱9)8}{�7t(&���BOj�=�zr���&����E����}����х|b�}�}�~�f\��x.4 �㶇�co�z�8��.�!���S�������E�:	m$x�Am�-�e�I�2���ӎ�ܨW̆Uّ49����4�ÝY��G掼�/n���s�JR�aq�0��:]2V/M�"Kˤ���ͽ��!���gz���Dt��ے^s ��a�#%`"({`�nv߂eJ0�����|��t���/n�*Un����=}T�$��e��=b_<_���^�|�&��ߒl���=C���(�2���2�n���mO0^���0e���l�&"娭v).�&Pr�b�F�̓�
6狧�e|Zm��zLʌ*<H"Rx��'�mA�8x�&���o�<�r�����x<�OR��P�fgrWZ�1(%#��?R��NΑ�v��5���b�u���$9��H�HWڊ�3���q��n�G��,M�:̕���m���&Ky��/��S�S�B��+<٬�G�v�"�gu�
�&�̼~C��d>���,D��� ��1�]|�S(��p])m��tGq����s�z%�%rq�VW����)N`R򋓙$�R't��e?�v������l�f�n������tl��ϭ9HP-�<#a�c��h�f*+��E�+<��'8�-�� �?�95��ry�N��)�G����x6A�*��y�+���̒�b�b].����Ϝ�� *im��̨��J�q��E���L�+~�H����. (�D�i@�|r�CQ�Z�.>�񌧴�Ծ|7(O\������]�C�e��1�R�&r�U�&�κ�f���'�8DB��.l��Z�C�8�B�<���a.p\�&>RǓGM�����uO m�l�US͍����B�w��}���e��=#���<�s��QOi��e�H�Qk�(.7�&��JP����Ό�+d�>�L�=�qeNJ���?�=�$�k����P,pQ�!��6�gl���2[��\�/��m�ӵ��9�$����<����&����>ܾ�p'݋�a�:�=^NPk��G!�j��<�7A@D�NV�-���A`��&޵���iv���9�$�Is��+�������2��g-QuC�A�sy-Ɉ��W�.����^SO�.{�y�)Q��F�������]�%ZK!�;Ҙ�dK�C��-o{�������߸'�����C�לЋ����Ct�F���=)�Y���<ޜ	8R ���{���#<�w$S�v�o�[�/��F��B��.��/�=�z:��||�����e���Z�Iq��A���`�g�\Vdh���n�
1�ׇ	q_�W@�
?��l���*^D�6�J%�Fh�^_�l�j��NT״��dm+�}+]�@w�r�L<�7*ׄ��1P�Z�T�g?*nIh�'���N�9��k�,%�Q�U����@z�:�����y+,g&��������?�%�����Ȇ (Ȼi1��uM�/qӄs�~Ɠ�G�*���+�hL��b������\�������5�c��Վy�h08^3�N5%/�;ƛbȅ�j��ɸ����e(k���� �)�C:����]�/j��bE�_������?���|�͇rU=���Z���gl���
�lr��S!�a+u-VLɐ���L�<RӶ3��rZ�F��FX��X�Dϱ�������/l�g�LFH�XF��eMҦ���+k�W�ݜ|��uwǾ?.U�p��
;��/��K���g�~�-PQU8M��2�I��5�?�/��B������]R��5�~��(W���|	���2ĕ���Զ�z���@���j�?{kt�O��u�+/(q�J�N�hg?OM�V�j�z�,Lt�=������b�}�Q�x2t�-o�b��(F,�xۜ�]�G~IOG��R�b���<�#R�eZQ<	5�Mi)G"]<R幻"8.	�[�/�{pt]�o�Л�(�C&�a�D3]v~)�o|gz#��Cv�K�䉓E�i`�}��Ï~R��vA�9ri,����@:�H�g{u��.%�ʷ44�	�<݊�T����l�Zҁ��� ��2;5l�}��A�{���ѯnndMmbs"���&�DZ� g���O��b��}����.<Ӣ�=�JY��:��UwO_�ެ����[d����5e��۸\Le`I�U;�yM��D��·A5���c��
�g�	>�HG����i�>��>4i����I@|�5L���{`���TF��!�Lr#�
�����w�9���ܼ@��ʾB�X�Ge��W"������bY�f�=/T� mO �J*x�\O��ېԖ�-�=\/����F@/�b]�q:T)3��ič�G�Lb��aT�~NJ�<��Pe�/E<�2�[s�� ��,��b�{�<���z=|���o�Oz*I��ҩ�N����~h�a�dc��p� �|�l���-��Cӷ�����N�_�<|�[t��������I���4�� �2��qA@]�d:K�E�qF�c����$TA�~N�M*F9Q��34�/G�Gx�|(���B!����Wa���Ak��4�g��'PF������z9�e��Y�! 8ieYMK��H����5Yh�)~��/I��E����K�
����z<:l�OF?Έ�ƝP3Q�y"#�X"~�li�� \��6�kRߌČ���iQ[�f��ݹ�N9a�l�k�&��+K�M��N�J��u��X�� �>��_[9V�m���(�o��FpM\>LxNP����4�����=e���4ț�M)/*u{Tye�[a���trѽ0C��mq�4m%2��d�!�Z��mU�M�ĕЀ��i}Rϫ�R"3%9��kd�M�V��S��zڃ�n�@�������n��;?Q"�,�h�F�nr`��q���Э7��\ߜ��ꒂ.X�)��b>�����
y��k�3ɛ}�<`I4�����D��#�u�W��Y�R����?S��W_�]Nu�i�&-�+h%4�:�����w�����������d��f���:�����g�[�wqҕk�rTK��禆���#BC���$��?��MU�n�j+�����ho���M�Һ6�eG_~O���18e�S�*�ԙ�0���+&��� ����ґ�4E�[K��.zb3�qW0���@���Mg���z�D��0��_�|�/-S�Tԭ��oB|�G��|�a���ub�����?�7����Y���x��)#U3��,{�`��>}_�!���:n�r����Y<�g��	��i ܊%�(��d%�,}M��q���������_l&^˼�7�)GbF���\_>`�:Rb�4t��J=m¼�,\�f��������m�U���?�]����ʁjo���Q�#oG$�uҋ�9�<i��{��Sےα��.$ܘP$��l��/���d���P�$ �jX׀ &��k�el���$O�q�f����bfi��,`;{�:FW<�و7GY���b޶�X�C!��Ł���"i��P�g�u�~��	֋`�
@9�m�;�N��q�K�}:!T�҄*!j_���[/��]4�>^NN-�9�
�Fr��p��K.Z$}���ip��ۆ�Qt;�@���'&��3J��RC�"�#����kV}���[�DS��`�����4��t�&k@�61��e��uu%�"�#5]�᪢!��=�.�r*�ĂRq	%�1-
������hn�}K��bl��������v�M��ެ��g>rƭQ |�'�4��*�n"�bJ3��`]���ԺB)bO����阢s�����t*������%r�E��!���cl�uߵ�*��!¨��}� {�F��{]޴:)�0�?���G79WU��v۵E�_6����CGb,��:��-����1�|�����s�����1)7�����[)�^(��������
��.��!@=�.r���Y�$b��P��,̷�]Oh	QJ�ea��wŉ�X�/E�8W:#ߵ>�3ytW�TK`��4�`�����
B����x%<`�5��s%Vڲ)A�� 5|R�/oX=�	�z0�ԩ�q���s����L2�����!�����I��Y?��t�l���:�띒Pm�� 0��(�G�{����zD��V|4�U��_ ���\��"]���2���S��C�+��Dj�M��}ϊ"��1��+ E��K�B�yy�n���^ ��o�\���@
e9�����d�tr��b��������������sl9k�a?h�F�b���	(�J*�\���ߠ�]5��L�;���a]��ֆ�7� �>K�A�;�
�5� �3�Dq���,���)�+���fC)���x���T���r%� �t�˩�WΦL���0�����n�S��5��8��w>��Wh�
����K�O�=���^�c�%���mY8���#��/�}]!d���)dUx<񻢾�_�?�Ї�E�j�HWX,y'�����@�2��BCŰ����q 3=Hα��YW���N��X�5�"2?S+;���26A�sfG��V��\�x�:��7QE}zexD��T{0�|�r"?�ի���(Yo�%���`��ȪM���N���G�i%|'�B�ˬ��4���xh//��;:��aq���Ҍ���Ō���������t�䬸#�Q����r��|3��l�Sw�O��8F�������Y 	Woc=����##y;�",KXO���O�"����禲բ�.�����J�G�/bQ
��7�s�k=;$$F���{���񊫫��4��r�i�1�|�����G�������(��#�5K>�;-�����3�O�|�pȝ:��� 3,"�[���Y`w�=�<�Nz�"h�3Wmg�o),�8�#a���ѻ�V�{�QK��HΎͽ�ǰ<�o����+ed�#{wCz6��kaK./~�k� M+�lT�����y~{M�3���(U2"� ~����~j>I9���bѤ�z����y7��T�����yA�k�KLY���$�+B�f���aR)�豿�D�ǐ-��G\��J�>Vh&|?��lt����AG����>���v>�]覈��W{����,�	�f����c8*���]��
�C<�-��j���.
��]k��܄�	�A[���|} ۤ'���4�O��M�h�K�WTy@ҤxY������-���6?ԓU�m�i��T�� �B�t�}����Vm[�bȚg�'�!�O�J
7���>h��LǈQ�MEZm�XH�&�''l���ZH5�G�5R�`H�u[m�/'���%�����cS�G&��!���j����5�z��Z}���~f����P�Q�?�r�£e�)w%�Xr��&o�ІpO3_��/l�i2�'�)܏��\��������({z�-�3�n�-���Y��ٙ<��U}x��o��.?�R8&LHB7FQ��'��3b��\f|F�n����L{����|uO2ǽq�Y�p���e���JQGo�DF����g��1�<����n	�_ݬ�gF����� �)��L,�j/|��krb�+��u/��C�t�Q1��;����?x��$�ԭ>` ���m��v�A����7)$�
�-˚�U��٦�r�yA�}vT�:�1f]�v����wx�K͜���M�n�}����Nf��CV6����r��Cm���bm8��0G��m�����b��,AC2��$�#P��Aᚘ���HyoG����ur��_��ѝa�|�2���lkR���8ۦ�ʘ��'�RS��+EX[)qjy�r��e��h.\)���7t�p�%4í�L��(��=��ܲ~=+(����n:�}����j��Ndv7�T��o3��:��7��,��A����Ǡ��4`OF�� i9��{{��r} #��s��I/��d��~�#h
5������A�m`P�b	>G���z�����<�-ZpC��}��&��f�$��,2��t����W�ݵ�#<�����6�2�H�}�K������;1�</�v}Z7��@�m�1�ߟ�'�W�P��__� �.: =l=�lx#E#<��S��:�i��BE�!\�U�ƪ���n^���'�_�1��J~�n������l~�`m����Y0.8��G�uzfL�W3�ȨD��)sF]���-q\$�FP�E��V�5J7�pՔ{E��J�"e�c��^#�^>��p;��y�����)7b��[��n�1^��m�=�wo�-��!ߞ��(�`�vxِHdn�"�7�4Tn�n,���m����ZM�����~��Ȋm	h����8I��*��#XU-�'�>S��C�T(QO	��L���][<�f���ݽb�b+fuq�:����R֯�_2����۰�Lw3܅����u ���D�t�m[��+���{��Oz�<u�N��Vp3"<��^�@8o�j�.Qt��,��F5<�FN�K<SU��P;���kݷZ��i�#�e-�L8�s�������3f�W���v=�U(��6px�}qO�/Kd����P���@��lkO�׷aFҵ:��3~3��� ��%�����.���}4���$޾BC���F�R-z��x�k�)��p��� &k�_S''���c��+?��6�< �Hr4m�DS����%X���9˄)�'^����X�[�y��bצ�c�2g�3GeI���A�
W-�&���/~�>`�\�T���W�T$�}jΩ���[�!���A�&u\C��j��de }��<%�uTc�n^8�۹8k�>�o.�oGΈr1�Ӹ�� Z0�)S-�̕�v0X��A����5���
�2d���D����;/	�$�����
Z���5v˄��7�sŵR!�ށ.�@t�d�����k�"��;���sa�h'���%�ĸ���,�p�n��d3��;$4���R|���&؅N������LAֳ]����5�;"Me&%���p��=���{���b� Z����1o�G��@$:4��,듵6,��K³}sG7�(d�C��oc�h1-2s
48Ժ�'�d���6!-�l-:�
%� `Rm��	8j�K���j��8(��S��)����`�>w����#`�E:gȄ��h[�C����}�nC&�Ѣg���\�kk��űe(�.�EL�3P��iD -�TKgj�F�H�d��(i����1t�����LfS��h,���q����|tV�ӵ/��#D!{��wi���k���}8�o>e=�����1��v��V"|m�}������!A���>�]D�'���J�����OKe��Y��1xW��#�[A�ӊ4���u�>p(��[%��7]��ata�[I�t������@���/ Xz���P�b���}l��Pz�%��� �|u�n�D�fK�?m�d�)4S��))Ი�E�t@��P�0z*�ăo�IEN���`�x2�a\]�	�T�e�_C,gU������!��5��ȣ�Ҝ���袟;��
��U���@�v������r��'�8@X'�ʉ�dkV���I�Im2c������A�0S�1��?ۡ:���z�	Dӯ|0k�3趓/�9�.��7�LL�f�X�S�˷Y,�����Nz�l��<
�KY�geMjB`�i�̸�g����O֛ؓ�㝶��D1XG,0j��%j5�ytP��U4��0`�7M�6V�r�
#��&�WO�/�ue7����M�ŐsJ�F���N��^^ӄr��$f|I�\5$Rn�z�T���|�$��N�?gEN��zD����h$k�?�v\3$:��Y���pJ�\��F���U7��ݙ����)��t����{��`їΉ\/��q�����K��7������ӷ�<�t�~����3�fZl�("[#.��4ʽB���M�g,o�B5e��sr�2����B�U%V�SS-'���b���͊_�·f�׎�2.��W�'���{�L�
�#[�'�_1��!������l��z��{�j"1����OjR^���o�N���Z�V�Y�be�Z�D���⩻�ϛ��~'}�Xt�r�`$q(�Hw�S�VM��I͎�{��Yv�y�0��]�ٰ�Gaa<� ��'�����7&� �3d�A��]�c
U�N[Ȯ���f)#K��B�5��'��3S~���X�U�u�y��Tx�x�k_M瀑�=2TjEr�_@���{���|t�!(�'���G�}�����o�G"�Z���'�JΜ	s�]�Q���[W�o��d5V>��_v-�@S{�'?� ��
��+�d����i>3}����i�!��~?/v��zM��3A��P'ǹώW��3�����)$f�MP�.S|7T��_�X�=SWN����jd��=~@�\&fZ;~;iu_Sg��+X�I��Wҗ�F��xR���Cu��
�2���8Uo'��������ʮ�4���+е_��7y���?�K��f{���̾�/ �k�_��ݲ��`R�\��l8���y��O�8���v�1�3(4�O2�8��tJ�ܽb��۰U��ѧ:�MZ�?�Z��s��.>���ތ*�:��	�.��aJ��^N*�_ ��bZ��i3�0������ �B�a}O�?�r�\�+�^��?E�w�+��5�^�7�()��s���Fd���^u�$��b{J�X���	�ؑ���e��&!������͢�8�����6+q�.�5(�>KᵉZ���ňk�I9���6���oU��b^L\g�.�# ��0�ٵnS���l�t����K8����l?�!��q���]���oOl �2���^�w��5����%�������+����v��[���R,�#<p�Y��A��g����E2?���*0`۠�I������񊶖h-��m�x^L�x�1��z�q����_�S��`'M��|���ߣ�����s�rƼp�γ l�!�]���!$B�	 ��x�{�+�>-4��uݺǋ>�Q�F%y(E߫��2&f�S��v4�󃲎�����}er\����P@7u9 RdWh{��}u����+�Qo�9��}�D�D^��϶*3��f9�݈��'����&�8�/6I��ϭ�S����U�P�5꤉Y��Ǿ���8C�wj�-U��H��DƏ�B@�¿0�!�� �꿚!����gaТ���}���&X���_���j�V֭���hͳ��1nN��@@*�:�6�N�I�>=��˘$�iB8�|�N�5Xm���Qp�����gG.�pO��KJ��F�Mk6�����>	�����ƫ�q!;5s"����q��k'�⤂�$�>�քYk�z�]o����u%G'5 �Bu{q(D).�y��<�V�B �7�e�v3�[�:�Jф��mZf]��r�Tk�5;�6�2V��o���o�a\��8�1o�>�
m�.O#�G���e��jN �NS�V�����ӄ&Gcњ��Qrƻ�2�۲��Y��f9�,l`˦dZ,?��-0�]���#z&�ռ~��:W#5_H��}�Vz���qw�����j@5������!c��n몐�S�)ۅJ�m�sTa�Fh�0���������>F�YB'��`���t�ܗ���y:2�������ELqh�ډ	�3�S���ߔ
������� P�τT�v�Y�D�b��4�M\U��W�X��0�����H��F�-�Б�״]-1��P�:���
5�0�(Q�ɩ�2v4|zwD}��rVD�Yy��
Pq�K��9��nKd����I_�sO:% ���x�=��T n����3�"k�`/aĨw8mV`�x]@	K�]Lb�$�(�<��	y�Ε�<���k����?��$�6`U�� �Xle{��&�N5��)BZ�=>n��+n+퉚�T�F�m��~(mo��4��)Go՗*��>n7َ;�*���wI�@C{�6i��K�U�a��_�ő��������Rl���9�#��g)0v_i��Qw����º�~�7�ǲj�����D�����NY���6�"hH�%�+�0`���6Ņ�~c�O�+��iFv�7��X6���"b��*�B6��a�#ID �����d��%�(��Kv�9B̮�wg����������z�e�o򄖍�>���m]l�n�Ch���s�i�7hC�lBbN���%���٬׫0��:"[�`R�d�T���/�-"�}[��O���R�[���zݺ�,6� �����Be&�L�
�g�扼#C�������>�ձ���2��Wtc��$�,h��n$��Ւ�;��0��u��8�f��咐���w�`pЈ�ڷ���w&c����U�q� �eu�¤�P�r��t2�w0y\.%"fg�Vz�,��'Bȑ�ӎ�J�yYȋي�*�����q@�h5�PP?3+��ً�n�� �����^�6�	��JК�ֆQl�}����dfg+���ؗU	�ܦ�Wh�v��`�����@�B�����Y���<T�Y�ҿ�p���c��娦��TI ��f�����4�`Da�6Q��7?Y�Ҷ�4|�ҎD���E���f�����R>Dq.�z`l^�bV�)�⪹hÅ�/�{�D�u�Qjz�\��I7'tY��~Y�Vҋ%����^�!X��#~�DM(l�����B�s��;�x�D:�����݃P�t��',��� ��G�j:n��5&:�1��ķ �1���69",<h�o�	�4�ڃq������O�i��[ЬR`�t�&Y2�B�KXUx���ܥT]����D����@j�vo�Y���?TZ�e��v������o���E���y�+<0NWW"�QE���b5r]Ǳ��$D�����x	��p��G������N#ڔܤ r�X\R�	���	���=��6y0!%�lVQ��<ֹc�z�	���P`|p�d���C%d�\G���sv�4��gZ��b̩��AQ�苝g4�ʭ��1�e(�v������|��\�;qผT�nӡՠr8�\��*̓��N+��b`�[��<�XY��Q�|'���Q�N�`8>��>�'��gKG��К�I�� =����� `��Q�m���� �|ߡ~���$D�I�^�+NH�E�U�dN,��Ts��e�;ի�������W�7s*7��_S�ap�ඥ����|��	;9=pO'�b\}����l_�X#S�bK���ʭ�i0��Oe��C�nM,Ż�gn;&�{4j��$-S~����Ѻ��
��ܨ�+T鳊����D	��juZ�u�{�4+���%���ad�X�Z��|�(����Zn6z(3������������Ǿ���e#O��B"Kgq��מ�����ά�4떇𞋗��-~��R�&����	u��'��\3lڱ�w!�5�Qlt�}��8QDc�����0�27���#��I�K�y��I�_߉�N�`&�W����ET�<�#J\������#�0��	@C��veܜ�9�}�	��euf���3�U6�S`�Z�S��a��@�z��/(�(oի����;�U���:vMF�L�9
������U�Zr���ڒ*��pe��E��I��論�څ��-�Mb���e��b4����Ր��X3J"�m��dl)��"*w(\���7qgK��ߐ1A���n,����<c�c�|��a�-�G��Ez�"�2���6G������ ����h�x;}�bx({�5���c�~�mdZm��N���N���B��ɟ��`�B����9����V����,�T�J2����̾;~���n��֖��܎�`ⱛE�C���3=Z���h!�@w�k�Z8�v�F+eM}�7�/P��?�}^H�����Cy���q�k�m�=T��1�{���x7�`k_�sJ���n��� 54���3l��-3h�ɟ�v�"��ı��ea�N�m�)1u��6�͉���]� ��C�1HfO�[ĘO�gA�4�\�=�i�$���⹭�ԛ|�rs�F���.���fh��8������眸R�諄�0��}o���i�q����5 ���Ӧ}۴�P�%^ư�%0q����eo�3u �"O�nIru����|]���d&0cK)L��A�k9��W��)��;2ϥ@a�5ݓ2(�d���s��;	�C����J�S��uAA��)����p[R+��K���?\ڠ�o��<T�SY6��ʫ$Ь62?n�5�b����Z���Y�¦�Џ���J
��k�U]F�1w��4v)'a��HW�P����e9��aZޝ��6G_A�zS1^D��ib�W�9���_J�q�:�\���G����Y1)�h�/VL���R��>]�f.�2�y=�;e'�U�~�/v�j ��SX�
;�}�܏Z�FMČ
]0���u���g Ye*8EPK3}�z�I�����̑�r!5�*ϒ~������B�/�����y�dA�'(��E�����N�7*��.��n<�g�^�u��%DGĺ����1���({�.�D�ۙdV��q?d � X��l��$� tޓ�w�|y����c84q���2��y�k|`��m"c�˰W�J�d!�2Q��]8���C�W�����tv1p��8��� j�U��oA��b�,,ۉE��%�[�H�׵m�y|��)�  בu�1�����O�r1�Z��m��ጙ�09wD߅Wk���nv�פ,���6�W�Ƞk��1U"Le�Dg����x�y�K��o�K(ho�)��G��F����������eT_��	4P&��<���k�`��ƴtd�@�f����35�g�T�x:�ݥ��!�TL� �O�!)^��?�'��v�0��cEd�AKfa[��ի��z��>��O²r�M����;��2tA!ք��5����_�<�L�Ky!�PD�\O���,�V�b(xB�c��jJ�&��:w��U����?l���H��uM G]]��ʜJpb1��/�RI���w;Acg���# <�i�|
��g��4�TWK�"��4՛��N�[j:�S�Z �-�}?��I^ur�ȣ�����~pu��h-�RHN�|Y� 1����B�
_@-W�o�q>4��_����� 1܊/�����g�O�_�F�@�A���%n:�h˴�U�#p-��*b�bN�R#|��U1��]�yympi�*�v}䂰ؠ~��CI�/�x������bp�J�^aj�T��'��3�����0�ی>g�3аl�w,X"d��딍��o���K^����Wl=(�J�5����8+���s���ܤ�R:e��3У>+�9`a���5����D"�]H�,��W@�0�Rw������$���|�|!�"��|@���9w�%�8�t���{3w��!g��Pc@�|�I#���\�������1H�� ?��?'�zp����y���="���+�Fg&D��I���J�4�{��vj��"sԴ2�&��ܠ�22��^�4���A#�R����{��#��KU���b��X��R�g���<�]���;-�u"R�y�3ʙnv&&���5̋*���A�H{�H�}I��;5?�+�C�p�oy��`@��\8T&��u�}bj?�L���4M�%�P
���*�P�N^�2�^��U�q���z��W�O9�;��`���.}��7^�7InO��������m�D��,���z5�鴣(7���
�f�|���r>��qA5���א7N�i`������[�Gw�h��PW��E�a�3!̸1��NS�!φ�b�W���ީ!��`��_��DLj/���Ln~���ގ��_��k)ڣ�嫪J�͆��2�l��n	�.s��S�a5�T䶺m�h����������2R:O2���tGC���D5����6w�:�BrLAO���LF�)�#�]�S�7.s	��tbr��5���==��L�D��6��X��y��.E['=�����D5pd�K��וp���~{����7mN��e6��Q��I��"���~�BH�{��6`!��v3~j� K��N<�^�^*M��z����a+L�,3�U/��K���XG(���-aʭr���t��x�'����'�q�-n�ln��hr��ȋ�K�6�9�-��x��}ocN��j���"��	��#��u�s;�[v�]�_�b��z��:�V�NU�[FN-�_�Y�I~�n<D��sA6 "�;��&�g4%���x[��8��iP��/w�6FK�~�
��eۭon��~l�x��Vy[-�86�Mժ��GJ�DJ�㞤��?��+������(�.�47�u��@ ��`����̽p,7d��kn~B]B�t�V�f�>F���ކ�朁啕VSf�����������0R?y�B%����r���XK��!��J�v����I�k�J�{H��>��k\r3�u�u��2n�TZ�q���N���p�c��#Rp���<g�(�$'A�}5�����vK겒�?�W�bQ=�O�0'ߝ,�c	��R֗�(�n$��m��&I��B��hcՎu�sX�bc�S8n]ؘ�Ѹ��7�<Ä��o?� �����w����pՌ�pz�
Ͻ�~9g��M���sx����rnF�)�ꃽ
���t/͹F�-�O)�ޑL�!�8q�KF�]��Ҹ�^�#�}����A�y�朞'L�ITH��,�dR�2�d�U֏��Ɠ��d����ޗ�∴f���EC��6��+\�k�	���tt!`5 K�A��MX|C��]=��|v�,UU���T��<��݆H4���׸*�
n��]f⤠�9+�_$�Q�a��N��������)�--��̛jkܾ���i-��}�pQ�'�	"a�*������9�f ��骟+ �#�����r�L���t^StӚ)6�N�#�ZK�L�6ƪ����o9�>�"��{#��������������q ��86$sih�7�$��#]�Ĩ��,~$4�����p
S05"���`�`*��u��IR�7�P�B?�����'r�գ����u��E��1�r��E\0��d��wß_�[��J8�5���9���L6� ೕT4!��9��GT�o]ڶ�^b�&��{`�(�D9d~p,C�l��������=u(f��RK���*�K��k��K��#,c���}W�O7|P���<�G�rgF,��
�:�5M�ͩ�`Q%�\���#�`�1?N^2��nX�F\��3u\TW���(���*�xOJ�T�������]�%�U��A3��=-H�U֕a\"\��!�
E/�(�}e��G�:��G	�����f�⹱ �(���xa������x$�ϙ+����47�Qb4A98����c^ѫ��d�ᴮ����6<�RRB�1V��(E/�r��Xn��/��t�/�r͟���z5!�&�Ń>�2�xa'qB��ԩ�r�t�;����q;ߪ�}q۔��DGp��~]"P��W�ñx�7!�L�DL�5/�����9�UQ�j�5���M4�����h��WS��[�Ww��*f[��f=���q��p��Ǐ*\v�d��H�Z�٬���7���\]��Q-�Ii���t�S���ı�l����=�I���i<��
A2֝�IhAx��I���C�o.�)���^d���K	�� ��_ݛ�*�gd7Oy�1�=��t*��Zu�@0?Ά6�j� O�fj�y�#�"��
6���\�G���\t ��
����"l�$�/�8�����3��<���DkP�\G.~��U6�D�K���F�9����=m:$���
�F���g��\�t�D01GFgj�E�g����S�hTO:���mb3�+~�$>#H�2��om��� Ϝ~-�2�p�gc����c4�9������Jԭo�/n?a�4D�+����豂�v��l
:{|C0C�0�����W����@�*խ)��c�d=��I2�?��0.��ܿW�sx�R^�������zx0��	�IE��K�N2q�YKg�$=}��������o�c�|�@�؂Kf��6V"o�Lsup��������F�B.���W�-u?���I�y�6�Xì�	�3o�#3e��Շ���宽�� o�xf�Ut9�w��ti���ja�
���s���ru�&�P�7m^���>p���:�4X^lh��r��e�L<����~k�e`4<W�0�� j�ӌ�q:`P��KFw��!��FRV�Us)���`⪛���Knm��M!G@�����2M}��%T�����NY���D�ٷ�'7�4&�lW��ŻP�8@q
�?I4�$�c�	��k"=G��lk�W$ߎ�@35F ʦ�z�����8%>|�4l�4�ʯ�؋�`n��l�D?��� �I% �H��n5�(Pd�"t�lHA��y&N�*p�0'��A��l� 4��("�'�V��s}Gku�RSY��]�,(ĉN��4�I��K�� /9*AmI�@c��L�!�G�E�A)�����&�.m���c���[��xs���j�G��-��N>E1�ݿ)s�ۛ����_��ޔl�7��١gX�&b>In�T��a��ql��g�&0��&��|��]��P��`����&�n�8S�Du�ߊ`�~��hM��/�Y�t�`�ե�/S�p�w�΁sF�%d ~��>� ��(�A�S2�7����rg=wV�A�¹8�;a_�bf����P�r�J_"1�Ta˽BN�К`����������b
׈���٨P���R���,
�f1S�:g��X��	����Q�r��������E\F�V��-��7\�I֩�-� �Z�6����Y8�3���#�+/�FY�{�t��
M���� Tɇ�y�ڃK����@.�!�S߅M�e�����;)��Op�p9=�C���݌JI���0쓣�6��>���X����Q�Gn.�%�́�j(�����Y��Ou���6؍EyHH�B�A���������@*�x���(=�4�8���]���W�6H~�Y���?v����']����
��I8o�0��Lg��Sk#FeR���#��F�����S��a����2߇!���[}�=�xIC6t<������/|?M�@\�=��j*��7白A������*j����c9�,ҭ�]�	P�h &f(n��j�8Ÿ8u�	R����#��Q��~,��@ Ƿ�Z7,fQ�`Β��NR.*���w)�2�@�E{�[M��5���6����8xc}��<��-=��-�s�����b��m|o����"���ʅ���W�7�U�N���ǭu!6�#��b
=8��jw���cI�<:D���\iL/-o��ɥ fIM�纎���_�1�o�����N露���[9V���F��m��A�w:y^^�C`/�0�~��[~c�{O�S�^�V�8Z%�<P�zI�)��&0�c���Բ�
�h bo�¾�ʕޣ����эe���ө��-���Ze���7��6B�v�F%c�sqf<|ah�b��%��5'{l>��p'��co���&U��}��S� 4,�3;QF�2C���3L# A���#h��A�(���+���(��q�Y|a'79Z-ߘ��qQ��?��1���k��|�";���Uz��= �&3����[�v8ܤ�*� xͽƣc����0e������E�?�~�10�3��uY_(�Z����+����o��7SSR-��6�ĥܖ�`���c=�]�m,U��窱��
_�-�,�7�vn�]�p��Nm���}��8����}@m'a��CD��A�ZEO���f���8��k��uRq��TK�i�=��g b����^��L��.^@��Oe�|(3k��VX�nU^����>+�����-��Y��biꜶ��ؽ��٦8]F����-��6c9��yRJ�Ķ��AP�1����w.I�*��}�N�B;W��pG�������=k�tD��l
?DQ�O�7Tz�W��� �*c��t���ԗy�r�4�d�T#�����x^[c`�:*��5�UM�U�:70sd:J�8���ٶ�B^� �L(Mf��� ��XB8E���Qޯt�9M/}-�(Ѓ���i-f��<ߝ�����m͗hܟ&J��G2.�����֒����p�N-�����^a�$mӋ���N5$���>�@��M�-�P-`�+ȎJ)���;/F��B���&@³{�!V➺~_>�����R�4��
=�ă"kK��\?@��y;�vlٳ�v���~Y�H�|�)���fR�����u|aɹx��	HH�$g��~V����ܚ�z �YZ\��c��`��5�袷��Ot�ȸ�EI���Q#��T:�� �}7|,�HW��iΑ�Z�:QBz�Ϩ��v�/NE�0�����,5�L+8�"-��'��r���UKb\!=��K���BS��o	L��pc߳bt���1����n"�e
��7����NP�7��44�Ϋ��ݪ������Nˍz>�\�E�&W(E7���
���~�J�O4[�D�I�Uj�A� �d��j��9�eA��l��(d�z$�?���C��A�]�,������7l�RnDi�Z�@�nK��)�5������ L��I�F��R!���F�6������.>���gw�v���]3w�D$9nS����ɨa�%H���t���=+5d-8݄�E�1)��b��D��>O����l@t����YT�f�':5����ր
L���ش���B Nv��&1�fbB��G ��;>��m�=�6L����≸~�%�/���M�|c���XG�7<�IlW�Ch�w���Z�;� B	�1P񭱠������4�����7R���j&�w�
�<x
;����>8�nߦ�G\��0������qkv���)PՊe%��#�����A���w�u��挬�V���Wl��IktR�U��a��M�7��Nĝ�r���5k��B���
��Ԧ����'�ƻ@������]�G�ܭ���>]\ �nz�uR��H�t�`P�����Y38�MQ�*�զi��=���%s�銌�)J��Y�!#�W�.V!�u�$}����l�e�>W��q �Bc���%7r�������6�mag�����'�����3�e���ɚ^J�/�0�A�rl�j�P��	Jb���j ��"�\���l�Rsm�dCf[8�1\5��Љ#�ܤA����&ҖX�ګ�`�*�
:�$}Z�7���|�6��m����g�$�?Ɏ�'��u��^��M%]=־9uM�*�&���K7Yi�;K�{�Fx7�RK�k����1�:%���[Lg=��S��=X#�o���c��Q��EP:��ej�g:�y��}KiS9��8o���Bu���6�n���b���������e��,k��A����q��oP_y'� �:��>�~u��aG}ǣ���"�����k�HH(��zSYT��m�;���t���������׷w���qț%K7B��D��s����'$�F�q߂j�@-��[��Pv�t������P8b`��<0���L.�3���R�jy_vU:6����#������~�z|�ϱ�PB�ixZ��RE\,������e�� E�z����NI����nˉGJ�ϡAA�ܪg���˭2�+Ѭt����p+�k�w��XΕ��d�v
yc*k��j�?@�+�X=FCՎ�؜'q㱿����n1�:\���fc2��0hJÐ�._Ԉ�<��	��NY4�� ��C���Xh���һ�%�<Ҕ��L�Cw�I�����dúԿ����|@������Ar���}�������Q���V�b(E=��L�p�$vYiӐ�D�����l/�T	���J�ב��9�=꾏���>{��8`NSRf��2���d.��4&腺��q��98�S�.V���$A�� ��ry?զ�!0K������&d�m	�d���p�Z�R�koS	6��;�u��	�"j�܋��~�ێf�+��~��v������]6�MOo�	v��[�Dg��\��/a���yU��3^�ZjO�J���v>e�,M�_�s��@�>ξpk�z�C@"x�ᅝ���e�\�Q�?�Q5
1���QgB
�����D���V�7\T����u{�Xhh0�*���{�R/�<�Bp�x�J�C�G�fUN۰�()cV�(�p��^jE*��z�f��*�ٌ{ޡ��^ke���?�|a��_4���Iv(W�#�^�
��R�%�Y2�INIl�4� ��x��Cb,	7jY�/(mpVl#7)�E<x�y.\�I���Jk؀ݻUi�،uR+q'ćPg��
�듮X'B�"��7|�+i�����2�Q��S��[���0��hr���c>{&Y�d�e�P|�Q;���f��_C;͕?t��j�<���V�q��<�(�V�����G��ʎw����8��Ի*��b�DN��V9�y�J��E��@~Y=�G�K�s�6��u/p��"=�&�����/L�u��6��\nrxul�\c����)V�'"�H���?�XkV���`Ɣ���耼��ńkK�L���h
R3��/�k��� w|6�wD$�ϣAPoJ��<�^��[I�l��[/3͡|��E��d��Z���M��w�`����;#��@{=X�a��ȧ�f�^å��81dA�� �:	<S����:s��	w���h{�H�9L=��&�qE��IF�ppIփ�Q	���Ao��M*�3�"�u��#�������9N��0��C�,
&(Dl���^��D�.����|Rgr��qd�!DH{c�� LE���Ţ���7��`�Z����c�e��tutl�C{*����?���Cb���f���� (7X��gL�pj�>G�C�2@�0�.���D1��+��5c�Y�-<���S�ߵ\��f}}}y4-g6�!	�����1�k�B�(�38� M�:���t�U�8s�j�pMfk͠PN���B�dWEf�I�������r���$^��L��h����S�_a�S]�iU�l�W��x���b~�4y'�{ r�"W�A>��֌ܐ*�9���W��(�}@|9����"9��zi��@#�:��p�e"IUQdq��L�7�NK�NXw�A��ؗ�ů���H��wr�-�8-�������[��{J�䋍#fa������!Y���g��f�Vq?L�?_�"��{2��A �͇Bκ!���o�(������Be����.�|���,`P��y��CfD��:0��bHNu������)p��ΰ}_��5fQԶ�ͤ�En7i��$<���K�T���4h�;��;]p����/Ӱ�����1��o�k#4�3h�.<E����r�ֹ�Ȼ��ѭ1��̇<A L 9���g������{�.i�BW?���!��L<)�b�^�㛤+H�D����=��C��h���R9U�(9̯=䳞�c�@֛;~3R� m�}����֝2��N�����\i�C��2�s�<~�'�����$�*9���^uж�oK��o���~�D��p>��p��`�� ��Z�ޕ��
��t�]�w�"��{�>�k�y�I�/�ϼ��j���s_��j�'F9���>����o���+|�+���d00K
� ��w�.���N���q�<�z�_�^�q:O�#�v��[j��k��';���5�!yJ�Ek���>'FH�0�F��>��T���fe�}<	KW����|� Ipq�k��g���7��%闖�AQ�'���iI�s$`u��0�ᱭ4��G�%��R�D��e��A?����vD��i�C�
L�����\��g<�����{c��(B��v��R��+Fws�
S��,���j\y�I�%J&��YZu��`[�I�� ��Mʷ��w��4�NJn�w/��7�@*�e��ᡌ9�"�1��l��р�Oi#��VD"�.�H�K��\Q�h}m0	�����H:J�Z)�WA�}�ebX��'��A��#�Y��JU�g?T�>��[�����z�㯐9��e+���i��H\=ͧy����^��Jq;��fm��Θvը%�"�Ԁ���.3�
v���jR"B>�ϧ�����C��_�a�l`�窝�Y�:@����-��^9�Õ/��TP���[eN�_!�=C_b�B�HA/ Thg �ړ�S�%��E��l����6U�(R�"X��0��k+�Pr>Gh_�eH��k�/l��AuQ���ޖ�۔�����&�Ԟ��з�lduS6��0Φ�pp�����g�u�%P���.��X�o0����낗��飙�4sK4��h�l��N�U��{����/h�i3�&M�#jT�c��N<0J��_���O�����Q7.C��&,M@���;�}�LFȻ
3���l�p�P$ۈ���7vr�)�z["��jc\�~���^~N�)�);	��V���sf(�y�m�¦�\�yj�l�(5���H��c肪i�U��Ͷ0����?_8 KB"�}�<��R�t����e�F�u��w�&G:�T���]��(>-� ���e���R�x������a��Rh�<�KH�pFR�3��p�+q�eiv�	h����G��D���שDH<4"�ms5��Q��qP��F����C^��h�e�6��D:��\���l���b�SuQWj��β���g����i.WB��������|�� ��jЯsL/�q�8�%&C�Ӑ��!0HW���<+��uK+�D!,|�u߽qI
�T�wz��
ū8���֞3�aK2	'oƱáڠ����Zt�P���%�q��e��c��p5U&�N/�b���tC/. �����:K�=F���?[�gG�N2��_*+�E���5DOB_[P�I�nn�$@М�����qXS�����"b~�ٷw�*�l�$�N�-U�&�ko���zJε�v��*oY�/f�nm��H̹P����+� �o�WL��#s� u5���X�f��1ݼ G�"�>�~|,�Ȱ��5��������(�2�}����+�j��q7�K�HS6�o^'5<�qA�ɢ�Ms~H�=^.���ѣסGÐ��ݩF+�S��s���l�)ЂS&�����+���V��'P����@�N]9%��T=�w�o�Pz0��e �������#��67.t�@��%3�eѱ��`��V��0OZ�� let��_~Be�k'Ѳ�@��Ƙd�,#:Ho��]�H! =}�;����(=	�]����'�w�P�Ul['����+ؕE�D�d�(I�g�67���d��,Y��!��K����[8~��\�_P��=R���4ަ��7��W[��
�ͺqS����ߐ&���6���:��4`���;��<MQ$4^n�hp̅�2����2(����Πdn:\���E�r��=�/M��-�J�-�8��A�}SWz�f�3�NgO9�5mە"ʫf_vv����*���������f�i�1X������r켾����z���u�-�K.�]��@ ,�mS�zb��|;J������?@ʶ鼧��_t-/.C��<'����e�ѭ�5
�� Ǜ�Z�����I"�y�XiGm�l]�/��@:���<�P oH*|֟����M�g`�jV�ԛ0Z�qrJu�?ɤ��"";"�G����A����\�Tw[z��u���t�%ҽ�D�~f}��V�;؏�I�(���(7rX�HEܘ�C*m�/�G����oB#�qlACx��M
lqi�0��ՠ���7�ݨ��G��o�_D��fL�pW�DS�9#5��w����]=��&:�z+v%L�g�����>Al��
�0�u��\�Yt:�2�T�A�Q��V�q;�o"�3�5p�Nl�g4��?)�w�ٗ?��$Gp-P�WF�_�c�FZE��U��r�
}��#��sޜ�l���}wXy�8��I��".x���yJ�)���a��w��oc8�M"��R��[O���閠�A�~�*5FXA�N�^�k���`(J��T����x���-C:�v���n##�3տ�}�����%�\�m�Zy=3	"c�o�a��b��p�F���Zm�e�$��۷�����H(���S6��+aޚl
P� u���:"�����J�(wEH��Y�J:#E����@�h9����k��TzD%J�nPS�L��;�c%읕��зjr�EKIc'5�y�mf|n���QQd���Ύ�"�#�F��7"le�gr&��ͬX�U!M�|�2�t����5�v�\�����\��J����/�n�*�
�rb�ג��iǶ����Gd 'ZSG���G�����V�=S�vV$sh�u��񈱒��1t2L�i�Ւ��reiywu;�%��<�;_�>����O��+�i�
� -\a����wajw9��Wqɪ���1��FkZ7�j��
�(X�ͭ7�W��q&V��a����:��Hu��C��9����Im	��C_�}&�lm�bTĵ�`eO&�\I1�����$LBw!mfT��J��=�Yh���1P�\�Ϝ��h@bZw3N�X�R$TK$sݝv��H>���7C�
e��Y@9:ȍh����.A�$B�6�3(��xn�'2�C���0~��t"�JR�`�;w������g&��n�����!�w�{X&�}m��'d%B�.xy�-~;����ͬ\
H��+B(�?NI|A�nu�_x������p'mЍ���4ΚA �E�T q�C�:��Jqá#ڼ!������l��.m$9�K,F5|o��w(9߉'Q0c�j�GNQ�4��C6/�*�hC'P��h��
���flq��4L�]�����j�C��"�!l!��!��c	a�YE�LJ�p�*Gn��~cXED�N��{a���5gL.�R ���Eڬ���8u;5#.~hi\�:�3�3��wuT'�0�ٺ��+"f��C�ØS���xI��Aܜ���&"���6ӫ�?C���;����bD��%ȉ�Y0-R��t��U�_<7[����r̟�3�	�&涒�R����P��~2��[��r���Z�C�h�5��M�H0�>��`b���������3�m��a���qi��Gk��t��!�G�O�AJxV?��,g�ͺ�9�;0�6ݥ�|�!J�VO�Jxz�A��?eE�� �.���M�V��sj�s�$��f����-���H����
�Ǡh���N�4Qv�}]URس�������_B�C�B]O����}����9����8ym'�b�i`~'<��~�D�3���{*���1}X�t���Ȭ��ھ���@��d�
��ĕ���~�;���/�e�?��,�����	�o�E�۶}"=M�1�W����=�GіF����r5-o�����P
xi����վ�����t�7n�z�"�(m�^�H�.���i#2����RmWK@�L)���n�,U�\�6ς4e :���׆^������䔖f����Z�.�Q�4ؾ��0~���6��q@��ᡠ��?|bь�I$�ي���L(��H�?F�8��k}�]�d����%I-���K�>v��>��f�+S��*��w*����
}���a�K��5��n6�r�6I�ݧ�3e~��;H.y���}��)Xݕ�u.~����k2b0�v�b��(<���k�
����I�J��ӽ�/r���Κ��0����9�/\}^����Z)�ոJ��\��mW-sI�NL��߬���ځb�O4�8�"k'���b�ǭ��ZY�dv�f�`��ؓ�^�r�c���?m�X钠�u0���/�Hu�xE#���:�n� }��v��i���}r/�^�g�ge��9�V=�&��An�/Œk����PMU�qJ/`����[�3�۰EE5�ꆪ�����j�-I��q�?ʋBN�7�����w��Еz��(�i"j O!65��M�oNZ�앥��t\����4�)����X��|�hjն���$�zo%}Fq��H�O>�Һ����ȺRe+t�x �8�r<4�o�N���4���i}V� �<���}D�[��TgňM�U���m�4�EP� ����SQ�9lbZ�L�ZQ|-�:	V�/��1�h���>�����Z㻱S�F���w��i`��x�1JzH���T���Tn4�e�.�п�t��~��5E�b�v��
��b]R��Xz�}�_D�iK�H(LC�p�`�;;�˱L��˦�:�B-�Ć�wxjIs� ����Z0����R�Z��|�Fz�X7$�r�t�QF�|��Q����-5L0����J�\K#����%���\j��\��]���^j�� �ͅ��ۓm[�o�>�q ��������@M�O^�bt)R��_�0bW�&�Y��GB���7��\g�;���(���Gz�k�$-57�u��id	�|���F+3AD��u624E1��beV��3ɑ�I ���6A���**1Y@�`��8�~�*�߱�eI
4qV9m6-�qu����}@�[��z���A�D@��K<BߖR�3�ZXԾ�pb�NC���|�<I?�h�6�ks��]�mz�G�	m��цmف��[�L����\��Ʃ'&A���Qy�9 �u5;Q���i��?Š��'�>t�`����������T{�L�
7����9y�]��#y4La���N�T���F\ց�Yy.�
��L8�v@�6);M>�Nd�ȳ�KN����MAE��8к�@�'b�#!�o���X��ۖ`3��=7��4�'wMy�$�Wҥ���`�t��b\�)�I�!n�6=���G!�m�;�XY��q�E�?�ֆ���{<�/��X �HwM^��Y�n� ��s7�	? K1� �_CT�x��b��#aK��F�N�p�;�j@�����r�ײa(���w�E��El�d��u�b�6����_%
-T���)�a��02̏�m�ů��Ɨ�zg�\��(S6Z(�z#iP��m��EH欿�좉yc�*�jl�,{ݞ~0dNS}�xY�)0��a'�uQ_��~���>,xFoD�uΠ�ڵ�:��DM�]PC�/%Е��ILL�&
&[��.'�B(	+Q�`�Q�e1b�HEL�?�T��A��7��2+ؼ�+A��/V�zG�~��u֤<����b��O2A�q;Y��]9�eV4Y� ���):%���;���������\!	?H�� ��?�N�	q��%�l`ݲ�|�4]��W���e��\ގA�ن���%X�m^>H�w���F�Qp� �d�.+��U����)�+8����nّ��ipYW�TD�g����8sD4L�'�݇��*����h�Őq�K�7-�j+9�U�D���Е����r��@C�b(���6w��=�6��EP��7V�������f���z�ܯ��h������ID��bT�Fԓ? yՄqԐ�����-�*�#��$3�L�ӗf����Ӻ�"c_[��w������=o���J ���W�Jx�U����G�l�`�*g��o�r�AO�4�W<�SWsD��&g��3�_���L頿�sƵUg!W�٣��w3A��Z��m����Y ������O4�ʦ4+B}����Y���t('�|������S�<&@��V�+���o\c]|�gHb��2n�F��K�6�[M:�&��� �0��x�P��F]@Z�'4��YOS��hB�3�6D����轫cW�m㕄*9z�i	٠��D��^xI�q�1;��sKv$�(���8�3Fu����1�<���f����ѡa~ p�
�&�|�	{Y�qB��	���J�&m���������ZcWc��߯c�i�X����M��󅨯%�b���m�_��� )l�	i�{ ���iH�=pq����0���Ȅ_��P��|�zsz9D�)�@ݻ�� ��z5�%�&�R�m��\H-.�+h0#��q�2{�a_C�v��K����l���V�R��BA��ky�|3�]�jf7�H�?��y|f�3*V�
k��9/v�@��7��@� �Yޖ���nuneC�����BB�Z1M�B0��i�j���m��jCw�l�9�)��],��u&M�c6D�O�JS�QI���c�Gϼi������Y�|�<�ѾO ��z���H�"��UI	�Sy�����Oi:�[��v������WVB.\�Ǧ�9P�5P�S��z�n�nؼ�$}|�����|L���%�~.}4�WG�o�}��O��40{B�S���?E��J(/�a~�n����	�t9����s�)�:��j3��g�Q�Ľ�/?�3��Pk!�����ٹ�����h���AV�ߣ�c�^W�"��T�ˋҪ�]YX�8K�3R��BS�߯WX��B�
~IhBԢ�x˧_q�%�,��k�����-P��ў.����n�"*�ߡ��h�7G$^EW;b����^������R6	&Q�v<�L7J�������2g>u�H���-~p{�jD�h�$j��ޔy��pz�(�5�l���Ĝŕ�v�3R\���O�cƋ���y�y�ف�#/��cT����f0�I\U6o}��0D���G�t�	KZ2 �r���>�?�a	�=d�V1bB�=!���QЗ�}�$�	9/>�=�u����E��E�	ۜ����*׉۶wuI��@ƫC��s���.~ŏ�r���$����duz0l�7�I�R�ߢ*�Er�	��,�d�0���c�P��l�y+׵��BЭ�'n�&��0�_>��n�wL[A�q��ĭ+d�t3<P�5)y�XP����*�
k�z�s��JOT��-^9M`�� M�b%z���0p���q���v�hd�6�Q�]�?b��ޜ�ݞ�� ���VK��W6ɴr��Mi��V$rN ��W���-����:Sn����^�QJ�n���1jiY�t�
�8��5Y�Id��f�M���%om�D�Z��3yy�d�<}Ԡ\���a�g/5�����dD��p@U��LL�Ԝ��X��TD]D����i!0ë|�2���DO�ŗEk��U���K�z��w�V7��N=��D���1�Wދvk�Hm'�Y0��NkC�����7��H�	��p�-
p���>�q�<+��
������wF�޲��s� /*<��{R�ht���`z8;��w��h�"{�l�m۬!�����\�s�����.�Ǵ���m�d�������8��<a�M%*K��%8��)�	@�G�����F�k9puU�0��I�c+�Ʊ�UsQ�4��)�פXS���������]�@������[�4m4z"�d���ഢytֳ���=e�9��z���Ś�_��Pw�w=��T`	���M�bioj��|�}�NcV�K�uTu F8��0욗A3���lR��,�H��D�����ԧ�����}ϒ�8ZM�O�4=ݛ�䗄x���tHV`C�5Gw"�E�E�E���\a��e�,�M��·���<�iK� $�i������n����$}Y����Rg���}���ߪ��L�q�xq��m����2�����/�0���rrX���0�b��oB�a>2;;��mf�B  ��0{6 e����HK��P�+�᲻�W9�[�gq.Y���յ��b���������O��q�����~�V�J���k�Au�XF�Mr(Wqc��E�?��s`�(���mn�f������p]Qa��)����)�KhS�1K8�s_�5#4|�b��-8>ф��P�Lf:Ow
���}������s���z���K�/i�C�_�%`}΃|�������Am)^`��.���a{��uEY�ĉ���x�`RJ���]� B�B��E����3NR(�P�*�̾z&pc� Nă·���<uH��\9��nO�V0�ܩ�j{l��IUɤ�F�i����9ܭ�F�	���N��Yh�2=�3$�-�n-jW�]��+�O���(KO��F5m�V�L��|e�9�%�Á{�1лGd�V�.GЮ�)4^���2���?�K-D� J.S�X�=�,$$>jF4((�j�`�}ig�g�Ӵm�����Bz�@9�YRs.�B%n�^�J�XL@ $P����c���/��FM/gʍE�c t��*�!)�^(�/b���U<�D
9{*�v�啛�+�kQ�ݨ�-��m�>�{r<��=���~[��6���!�)��B6��z�[�5�#�*y�HL�~v�v\\��t�<��b��e��K�sP=8h���-鼢��|��یX|��U��Z"-��pkT h߾+<f%=J����V��T>5�J  %��t.
GU�(��%���&��>�C��I����ɍ+~_C ���]����j��B����gA����1�k�z�?b��yE�&+e�{�)4T>	�#����lQ�椽H��9�FG����W���:�ά�w�d	����kr-@���ꀪ{7t��۰!8SA�2?�C�U}֙�_V.���/�ߘb�b���e�9��%��U�J@e�z�Tf�nG���>a�L�fZԷPZ���������%��\�񰉴��q.c�y�T���(	2�{���M<���_�(������qJ�N��7$-|��ܓ۝R-�_���~�?�b���Q�Y���̋��sbk[]ϋC��7��H�7i���@�����X�&���V^>��'(����Ȇ!uCEG�g�)W5�D���`"*ʳ��aU`_�Tr=m��|T��FaX�jy�x�HX����r���G⶜�����`r��U�1���^;K��l�1��YU唤G����h�G���
|�b��� ���\/!��-f�p_�$�*[�d��U�ɡ:��d�D�Dc���D�3�l6Z�j+̷�gH�<O:�������H�,&�1�������!�h�`�f'�?y�����,	��	�~�#���"����Kv5ڐ>��G�jY�	~�߬�������9�Uv�C�hS����U|�&g�TYrS0�������Uǭ������ج9���x���zi(�a~�t����Nc��Ҡ�wЉũ���_�+t�i�&����MC�+�CDxpv���#��ցm�!a�b�(M��d<B�ֱ8�Z�#����n4�k�c��P�9!o7�o�S�96��}mK�yXE���S7,�+j�d7))���˹�ލ��Ou7 6$���Q��cu��10U?_u�:�$�>�Dp��
Ɲ����D'������ஒ:.46߬H�l�	�?��w3"I �]�s�h�mۍ�����0h�p-KY����HG�F$��<��[�N0C�a�с �z�r�^�0P��]@KX�q(.�C��v�	��>Y����TA=������G8o�jvZX1�қ9m����S =i.�;��P�@�/ b�!OX���?Z�͘��:��"*ǰ-
��׼c.,B1,!�Hfs!���9�`Ԧ�!=�D;x����[}\.$Qc6=2Ѿ��)����?p/��C�*޴˙��FFY7�sb�F}�	�2�W���ɏGm�����됊@#������.B�F�<l���]�u����K�22&�VY�'��G`ڛ!��O:�������zS�jw�F�g&�7=����㿡4'�0Xh�i󂇛ԹkW}F��#
]G����`���NB��]�΢x�<l#+�YM/*�XO ��\$������-�i���������tY�U}�HuW.qչX �_D8F%%1�W�c_�>� �P��߷�o>��W�	�=�D
�*Z XH`&��ƺ�te�T��U�60Ȅ�dπ�Zv�hq�^;)"� �<߹��Y�`�;ū�Yڙ�:��cw#���sfǢ��G�pIw<b����� ��4��M/"L���nu�O<�����v{��2Oe8 Jv`�F��&�E�'{����¨��V��ӷ�(��}��9��1�e�c�EWr?̠',)XK�1��a�>޻�H+ ��Wf�E<��(��,i�k�t�FU1Y�t��+�v�՗M�"_պ-Ai�9���H}���Jnؖ��Q��q�y2Fz�~�G���[id��R�ۉ���.�8*��|�,�! E���ש�8T��.��O ��1�b����z@��'�ô�*�%��b�%Pa�벻�����srf�j�s�C'�-��ԞK���9�����N~�M���<�4�� d�w��X�6!9Kk�b4(��6.mh�O�vC�`f�����1?�`bķC�mPT��J`�h�\�y^��5�ڞ��!�3_颛r_�����/�b� ��D�MW�;�
��Pq/Zw�E��ґ��Y��������*P*��ֹq"�T]x�A��Ƭ������7�=��S���0
hW��;�$��t�%��)��W�_(P�h����H����ǳ�%�~��R8M���k���� ���N�dg�(�X�hsD6(A�G5H���I0fjvi�$8�Iqו�UB�P�[���)����	$ۖ�Q�t9VH���m���9Z����z���דBc���2)d����0n���p@��^�`}y)��iYhED_���q�PBj|��F��v�m�,��k�E� �ʅ���9�vt���e��[���'p��6� x��]]Y<�v/�P�`3�w�� ��.���V��R�>���2���.Bw~�����*�yYF��@�=���P��P�3n�s)��]�����L'����Z��FzpŚl'̆�p��DUsR��)ά{�9G/�s%�A�����)�}�����ؔ�!;@M�_�d���5�=Ϟ=�~v��\P��Ǯ�ˈ�Da�����d�����[�$_p�h�1G�,ޫ���y���-I�d_	P��k�&��k+��KAnDk��\Lȵ�|����|w~f�X�?�p��K��P��N����E�*��� S����`����5�o��.�0�&� l1
�_m��e�
b̧s��]��73+�&c���
K�V�y�R�S����sU����f�����i����ru�H�|�q�P������A���E|��i��h�i�ԃ^~��ͩ��ʼ�o"�;�,G-�ڇP.5W��d�?2BZ�S��;�*?��*x0~q?Yq�X���� V}Y0g����):����#�#��l���r
0��V��=�TJo�?4�B#/���y�Dt۱4¢�\?��1����{����v���4��d�S���������?�WG����Ǖ��1-1���aX���֨_�K9k��'4���'��l��UJ&t	D�.n���5�m{!���Yi�r�eC������P�����J_���/�g���!T���s���Ф-'W9�>:��Y	K
�s7�EP� q�w����V����fv�F��#	F�cIoZb`�q�j�kG���쓳B��	�]dlؐ"��[-R�q�H��Y��Te���k?�8}��0/���J(Tq�3<�d4��K��B��V׈�u���Ϋ��1��o �mE"��% ���i=Q(c��rƋ�pf��i#�"(�����j3Ր����w��i>��\���q�dg���Ptc�S�|{�I�S�iAԇc�<j2l�I��8���_f�r0֮�!��p�B`Z�+�X�#z�O�M{I�[�R2%�Q�o�*����"
R�N��R-�-  �R��A?h%(G��$���W#ѧ9)=�J։��� ���@2�B�?���{T�,/t�Hp�ؓ�rC,��̖�_��W�<��@:K�X�^���3f��;S5q���ƺ�q��n6��1t����D�'��n�Z���-��G�����I.ط/�1n\gk��$��Y���6ʖp�fX���ܳ际w�?�@j?2eкA1��8��#���Y]�`w�N���S��-B[�%�^�����5I�o��bC �XلGUx���U�q���n:f�^H�t�sȝ��񲶝٥+���
l�3�\�E�cr_ F�����׈����U�IkbI��~l���w�"����r���ӥ4��u�|�����24{�!Q��\{�ܿ0�ͫ9��7zv�+>7�O.�?��:+s����~x<�u��_m����	/�m3i}�C��j@6��:��K���]cT�5q�*�3io�>T�����43�1Ʊ�rD&�X(�.˲�x��� ����[M�}���<�j������`ܸHM����B�vCȼ#%X�=�f*�`u�k��&�-�$c߯R=��$\�P
��0�׷
r��S����k�t�U�o���ʡ��(�"p��D�|]g�X_��ey��#>T"�������Xj�9 6E���TJ�Vf`
�n_W�pF��|��@�:=�ֺ����x�ǚ1<���}��?���5�A2�8�.�z��[<0�)�R	&�`ƊʁBe����J7X���r)�1��^{·`s \[��H�����WBz���D�D}�
 9K���>�ۢe2�eZ�	&sK�R'z��×�k�N�2Y�>
S'��e��2�h/;�C�߽`�s�6�(��$�_v���9�D�5R����R-�(�`��ҵ���n�"�(�LC�҈���`R�������5������:/�����Q��9�����:S�GE�S��5�kW��c�s��3=�1�ʦC��f�C�xf�`Z[��t]�i�T�\i�3m��@Yu[M��W�Ʃ�^I:�gq���UI�k4�5*Q��<9%'w��>��]w�1|�|������J�k�s7�l�J��a�t�mTd��-���)���_X#��:p���&u�0b� �D�؄-��"�45Ne�D�Ii@gmY�_�,#_���V�PXZ粬&(�Z�Xl�%��'?����Q,��ס���SW^���ܮ��hU�v��R>�'`��@%
�b����uB��Rt�[�$Z��ٝsIt���T�[&�1�]��Zmf9��-�_)ag`5�����J����&�⯘�C0H��e/4a}*zA��3Y��M?�I-�(�r�>�f�*��Ԏw>�}E����0���!�-�&�D�˛}yy2n���^g�4WM@�'��K����Ӕ�k���5�=��%밂�jue�rYX�h��$�P��yF�"|Q�UZ0���5�F�-���H�:TjX;��c��Γ�E@Dq�4���`oa
^\�!\�?�ft+8��|��Mo�#�9�O�9U���FX.���g�NN��xI���!$���Ɩ����rҥ4��������*��w� �m�Mn��Ɗ(����ͥ˛	4�Hgmt*U%����m�����e�ǐ�s��w�-/�K.�g����ְ����$x��E�����;�,k>ݹ����e1��/�u�6�Ɂ�V<��Q��tHkoE3@<�.T������1U�L�w�� s�҇���@4��i�])�=��[�Әz����ƚ�Qk%eZ�����+H��H��:i��E"M�p�n�-�
7J&�7b��2�{R�RW���!=�e���'=,����Q��4���i�ןS<W[��/
]�98����K���P�Vţ���ǥQtP@�P��W��G�_��k��o5
ҧ��*��̗�I^�������������O4��f�l�� ���$8�DG��q(������2C��
Y�B�B�$b^:�W��
��t�PL-�ځ;��P����������ڋ�/~�Gvl��T�2I.��d4n�|I+Y�a�4��3�N��I�<�����=��d|����j���lr�pS�����9��7h�Ȃ�=�Ԝ��-��h8������G0������Y�2�^N��ޒ�����'8�ht���Y��I���ͻۆ��I�t���;�:�*��xQwdF��*�{�(K����M�aI�Q;�Ա9��f%p.l�go�m��M��b�l�b�UM2u��MME�{�J��7%��G��5CR ʇ��K��gM.0P���hR�zR^�F���b���NI��l�a=�%Y(��[Ĩ���%�+�y�^]�.2g�s���oҶN��u� �̭�v�Ă#N��H\�g��2yo�B��z�.�`�d�~�3��b���wV��p}��[�����[�>uYA	�W�N_�.���$:dj�:ma��_(M�����G	<��7(�ug��af78���-��l3mj?�'R˄�).��z/\O��W�	EG��ڏI�hX�H��'uQYU_��p�#���Y-:<eu�Sc������e��ǟ���[�o@=���w�o���FJ���$���o���j@eWwh��VS���HB�����m���5� �?譗���O�֜^�Б�y�qr�9�FD�7[���:!h�{(�d��� z������p�i�~�C�t�'�2	}��>7ʦ�������ל�^��E��9Q�Rğ��d�@�U+'��EH_�q�.��<�&aNV�*p�4&�}G���|�F�8md�|�S(:4_������~����'#Ä����s�/��gqPCj�A�� ��T����0t̳HD�
[�-�����7�l�:qaipb�������{\�17�D���C�TQSZ�D�̕�{�P4���̹���8�J�Tu
I3�o�l��EU�9����rd�2�<��h�2[���K��qT�l�2�0T�6` }Yk���Z�tR�����/he��g��Z���7��Qgě�G� =�p�	j8'�#g����ˮ�N��q���YS6Z��⫉��D�Pӳf���w%��7���d�-�eD�]����A+n�/�v�N�HwB��s"�+Ft#%��F*�����,��"��LѽvpD����3���5��(lۏz�`p��Bz�)Ĵ�JRK,�H�g�uY9IǞq�UuX���Zoq;���gG\t7��H����_q���`_�����&/�e5Y��\�Y�=��s�PK���Wd�����(A�
�����\.�z���T��9m���؀h�բ�y�s��w�Ҥؤ%����Ɉ,4�a|,4c(��_��7+�_E������^��p_���!b�1�ޕ��	AzWv�V�I�T� �xr62���,����/�K�}-0�rYRjS��t.��g��{��Q��c���PZ��{�u|n��:QJv�5VmE�"Z�����T�E�-�#����n���إ�W_��A�;�dgUN�3{���R.�앣!:�n�3�'ԏ�5�9�\-WmIXՋ�
8'߉ܗ�c�v�\��C(�ax�h����ݥnM2����/�5G�NF
���u;�$��I£#��P�@�M89�%���%Gw���E� ��m�Ц�겿O��jC&)���>��������R����˽eN��,�(@ ;�q6����7��*��9����<C���n�4"U@��b��^ڻ�@�u����9�o���2J���-k��Ȣ�ދ9�=��E�m�c�R�;
_uBU��;#�+�36T�Dy��չr�bL���W��p�M�j����W�¢�oK��8��!X�W�9����a���h >�����д�u�\2�����!n��ց����򬧤��V�k��iV�%ί��^-�E�i4��x�s�����\�~o��f��mb�g�X�cG}�8�eqs?�F�5�����e��S�0>]��aU!4m0���
�*2��g�h����Yǜ�|z&>���e��hXn��7�c2��������a��]�;��/�� JW��i淨����b;��U^�Ϯ�ӪVطʰG����Y�(u�S�ňXOӤTL����ޟ��	�J��|\�[�����bϲ1�0e�:r����o�@�U��ql�}������.�d2�#}�?܇ⳳ%
��g�\�d����Jė����cه�T�/q����,��C��8�`e	l@-���=J�'�?G���Wv�MB㔷|R>��J�K���{�l9n�_�qEt7���:֛	����YM �/��;���Z�Ж���h����V�8B�Έ?��(��nIx�5���J��Nא�aE��Ȋ�^>�|Ϭ5 ���Xa%���#mmE���� !޺�=A�Ԁ ���&��2
5yZ�U�~4����/���qH[g7�?+�rF�����L�j���	H7Rq�`}w8�����HM"iW�{�����R!4e��x�~��mM1-�p)$�Ҭ�P�t���v��U��&߲���5�d	L���0���:q��U���tۘR�IS�ߐ��M�uýS/�^�	���)�Q�&�b:�)�oA�X����GF�M�$e��i��$���I N��g�*� ^mI���)�Xf0��¬����]��W��E@��@��[Bw����xK\sm?:�sٹ��0$�����:��P�EQ�c�D}��L��l6�
R:6�g���G�L�1ѯz7\���H�Dx�I�����IpF��v�|V��d�F���-V��C���^�j��H�y�X�e	�E4��`��iH��}l_ښO+s��3�tZ�oz�
�H�sIׄ�m��y����
�2V\~O���jjf���)�ҟ!��N��#b�� �1R�g��gAkNfobM����kr�2QKXR� �״�X���e�%�M��+�3��X��C^~��Jv���m4/n3 �A||�O�h��C��s ؃��8�1�ҫ_��	����l�=��+�F��1�� �$��NG H*�����y��m��
��55�����vrx
p�F�a^䟂'q����b�3�LT��@�O"�#�Ea��0U	���9VٯҮ��{ֶ(X���]���x��[<��ks7O9�h�}Ƨ�n5�6�qE�c>-b'����	W ���@� �L<Rڬ\�z��M��#��gc�Z�3q��<%��U&I��x�4#���x��'z��[�dKؗ~mB����ΉF���}�ݒ--�T*��|#���0.�P̏�Нz	�\��g���&ýJ��h	�!��G@ґ��^"k�����m�5�h$�Sᆊ<Nt�mIo�V��o����w��nԟUxPb�i����h�o�@�I���� .O�_�n��:{Y��I��4[�#6?��e���!|�µ��4�{h���R�����ٴ�#���]!���jҧ�N������pravZ�Ɖ$��V���ԉ��Eb�t�E_�J���oG_��Mn��'��i�©Mz3�JnOԊՕy�1�y,���,�(g�<T�Ѕ�,����`�M��@s�o��{7��F��7,1�����S�@E.�w\[�$-G�?c�p�b/���cj�ۍ��o�`W�X@�P���{r(R�8ѐ7J��2�GQ^����򄓸?lQ@���f4,�c�I���r������I��{W]Ʃ�h6���SF�6���`�&�h0�*�n�[���a˰�)��ؿԋ%�Cw9����u忡��I=�<�1��Y��S>�}�C�����j&0���A�zo���!�M�⍝I�u&����5F픗Ho��]է8Rᩉ����������˩������o��u����V䭋�O֨�%��
�q�b�j%	L�lIK��*&k�x`R0�(���FD&y0�u��3��sB�P����Sn��İ�L���rGlr�{A�z��$����6�3ϑ=��r�p���+��L)o&S���vD��*p����@t�N���o���贈P��;)J*�I��9d1!�*@:f�� ��ת��i��/Z�o5�8K�SBd�ep�b ��R׉Gk�y���'r�G��w���5u^�+�A�J��Q]Q�b�� �) �Y�)�ڟ�`-Z&����-^Bݧ7����'�gxA�ȡCxhQHYg���A|�.�O/��1�܀�b�c]6[01��*���i���(bBF��r�lLӥ�ȣ_�e�R�s���%OZ6';O��5Et$����e*�
y-���xB�H�ocv��B|Ar�TsW��_	h�`4��<�j��jl�,�bd�tq3�e�񜧭����I�FM�$�����l�*8Wm�mQi�?=g��H�6uZް��:(J��La�1������$�իKo�P�$5��d�$���\OQ�L2�z#Q6���e7�VH�Ui�n�1��{O ��;h�"9����.3n��Y،w��Y���^�`f�5����?�i9��
5-i%h�Ԗ���t� �ϫ���	A��XBW��M��%=77�ϩ�|ED\��c{������������#>�$Dt�����i"��B�P+&��gO��D,�-_t�ɒ@�Q�>n�G���(�tr��r2I:��R$���^��fX�0W���gF�nm��i��"����٩�/��H2t׭��u�iH�Ȩ
��4�ltC[����8�[���DJ����8zF��#E�`������T�k��i`�G�pW�S3��c;H��~�a	҇�A ���P-��L~6�=�1�sYR���z#�|����Y�ӢBĮ�.Ҍ� �}ش �j>(V7���3���Ѳ@{�Q��
@�x��E@�k�}_��CB�W K�_�z��b���� y��M"����0؜%�ҟ��N���EF���ֻ�x�]o�XE�_:0E^~��$�GԑFe�*˜u�i� ��6R�\��a���=y!cn3R%�?�����>�����53a�åI ���9D�P�N$�4��0��*�����j���%"}��o�Rrt%"6�ڔᔦq:N�
���. ğ��X=��x%I�X|*��	xd=0w2�A�{b�'�]|h�&Wî�$HA�!���C�lz{08MM^�GiΓE�G.k�-�6\<��JҸ�T������()HV}����-�g�����b[�9P,�Ռ�3�����wa�Aj�)Yz����#,��e*?5�B�q����n6��:;�4$�Z����z��k��͟�}�X�J�F4��ŝ�:αQ����N!�lݬk��TnBO�^`�̛�>I��KK"���>+�mK[�`>b!���Җ�"�8]l��|�<M�l&��v���Ҷ���$�:���c.=>]�6�R�#o��@=[.�>�k䄸��ȓ[�F����H,kF�1/L�J����u`M�d����K�J5-����5
^��C��t���l�mf���G��hT%��ߒt�yY��hI�\�m�4�ʖpd��,��?���\u��/��%��G jB��	8D�m��*�ƃڜ�TN�`'GFՎ쵢�L����}��j�	�μ6��F���tYi��	�m=6`&ςS&��M��>c�eǙ�a��sS�$���WE��m�f���Y%�o�P�����g�v��`?��f$���XNc�,௟��zx2A��܅���e�g,�?��{��yUy���3�-ʙ��?�Z&0�*j������O�V�Ε�;f� 
�JO�Tz ��5��;u��L���U�X���u��t�U �;�����߆|>�qF}���W�ڏ��9�x3#h�^�F���3:2=?����d	4�X��� �?���_��7��.�ua�_슋�m�g�9ݚ�F{�_i��#w~���U�/
�V����S��PD�Ϟ���W��B���dn}�B�vv��{9R�<���Cѐ��w�F�x켴B��"�6��9���> �������'kpP�;��`��#�N��߬ɇ��;[bK1n��sh��˕7T�&���L���`-O�����\�^�J����f�[�1�
=#��3����j+���T"��o /U(��	�S�������V��	MO�e%�$���3j:t�0V��8@GH��a�L�j)|���P Vp�6�S9N�#����[�Enma�Jmj>C?��}!�X7����狑����&���-�!����H'Bg�j�d/Y� ��.]�^��fߨ�g `�k�P�pپg{��A�]�23Nb��N/�ٙ�	͓q�������H�C����G�3�sR��vmB?K��b)�zq�y�v�a,�����V���@Ӡ8�3�tAz���gs�Wi��8opg��ǔFX�*d�M1�_/���.�!8�]__$�*!��SXl����j1P�kDBH$8ޕJ���k�(5b��||���q˧BK�_'p���m�>5&�Ya�*&(�\��{��s}D~.∛/�&�*b1\�J���S�����4�"FԜ��Q�L��@�pY�� ��-r�|43ò�9C�=}��F�,{H9=u�̙�g��o�oh��e�'h�|�\��T?f�e��ڮ�-�(H��&���<���ac@�Pj�g���qG���Uܦ�R���؎���bl��}/�-�((E�:9��c��[iu~`��Q�dp�!�!Բ�͢+����ܢHM�~��y*SC�
5�>���f
`j|�5��� !"���,�����~�����:�M��E �x�Jj_*fO�i�ó�D����A4�d���*�!0x��� c���!@r	�N\4$
�nޓXzbo��=�ѧN#"I���](��@�U@汪/)-�e<=��g����m���V9f��WMQi��
Ql� 9�}A��Y+*Ν�s¹1���E}Zd_j*:��6}�'D����H<ע�v� <�C�i���u�Y���@��[�Z�ުv�m���fG�<!}K��)*A�->�|dL>(?�@�%x���®��sL`�>LOxS-�㖝�ߏ���K:���5�A[#m�P��!���+6Q�4U�ذ�Fm-x��l�_�!��6p�%[�Ew��o���l�}=�ҧ�oĭH�"2ˡC���x�Vv�v�o�]�k�� �X
f�ti`מ�Ӟ���%O�yW�9��B��%���'7ӓ'�������hy���tk��$	t����^룽�DO3�M2O=�
k?6�pQ���?٘N���5��)
X�d��u�Z=�#��I��4_��T���ƚg�����T�>��^#�duCN��"��J)��p+�ŭ6�E���)�Ws�yZz�q��L�8J��A�<*���
��k�<�Z;��#�����e�;%'�8묻��T�P_ͻ�:@C(�=�T�W�ni�'��j�=��]Z�9���8��4��`�ȓ7���SMށ�RU'�yB��'GL�lI������5>��q�1���*�_nga��!ˣR��C:)����D��g6�䅚�))�Ly���XHn�ЩZG�U��8�� �)ٛ}���c���6͆��^��1W>E� V,���ȋm.8hI���ƾ���(��$����H�hj��/a^>9�J�L�N���ʋ��kZ`�  4�;=�>�;="�@�!�b�}0]�N�;����8�MϚ�_\�A��P��K���[���t��Mbq��ʆ�!����ݚ�x�����I���w��c��Jj�a�)�y���Z�oc���\¿�ל�f�H��U>\�����X�r�Q�J~�.�T�0i��,R��1n�p�������>VΜ��tM�}������#�.O�/�@��Z��f��� �2�c%;Z�Ý�e�6�&Y(��[X����|V�)p���Wδ��������҆��QTE��)?�j
�k{���%��T�y�NyRB��ʈm�0�>�n{�)���#��4�U�1��[ �*���_\��T�KP�Cu�n���������כq�r_�EV�c�]��=��8�^���t�)C#��;nP�����`;v�i�>���T�l^0�0~3�Jt���
(�rj��̲���=Ơȸk��ڥM:�;)fsv�>�J �~q��t[�@W)�U��J��&y6�?����=�ԣ8�㘔�6����D4n��_jT/$?Z�Y}ޑ�)YWx~��{|i�*Hm:D�I�1���K�������q� h�\B�o�fM������t�Ǫ|��Wb�}�>�4ͬ2�-
mn�F�#t��$j�^|+�NQ�=/�	�Vs��ʭ�2���m�c<�)Q9�2l�������� +&Ng�М��SǓ[�"AXy�k����k����>u��TFR���>�p �<��A�7α��>g�,͟��"�����].Hl�z���e�t���0ȋ������/I4����*� �8�0�f
|���0��	ny���0P]�D�T�Ѽ����u�h׃��I��Zvy��۱VI�}}46��b�!�+\���Qi&ě9�э8kT�x��~�A�a*M)��l	��ͤ��(�l~b6�H�l���5����+�fxR��1M��dP�86Oy��g4g�d~4�Q���)9ѥF��ǚ�+]7t��Џ�膔!�"�4~6)(����'лʱy'2N�X
`fvM��k�՚��ݙ1�w�c�;��#�E�P�O�u�CŰ�;�.am����k�]�AVU���Ո0�x���i��Y�cc|M��
xѻ��D�`B�����D�l�H7��4빋א��'��5u!��B�2+et馠�@5�#��ώ��$�&ޗ=,/�gˬZ�,�W�ڞC��T� E
���C�V�9VI_�~6g�{���Ъ�1��;�;'0��22«��N�zY}�>|��E���H�hlUv�f6�m�@�:mڳА�2-�O�=����1�i�i,�M�/ｫ��R�}�����[W�Z���_��(Z`@H�=.�7!չ1ʰ���Syͫ=�(��Wޙ��f�-B�d�!+���/��@�}/�WJ�iUZ��/R	x�ԓO3���_L�H>��� S��������E��Ƥ�$C��a�n6:t�L�+�6��,\��q �ֻ��h����j�d����E�����31j%�p�����4.7N��"Z�e���!�q�\�}�!]������XC���ـ¶����2�<'e�e��<�<rQ2N�P&���{��$Ͽځ�#��{����p�l`H@
�y�M,([���>=��Y���r�`�,T�o�TO�fgQ�C#���ڻ7	<D{�f�~����[&�/^;w��"�I��k��-]>�Y����j୾�Z����{n�	1̌7��-��ѭj���)-Ǝ�2Vp��#lǳk5�u�ݟ�l�Z�R"����3���O��a��+��K8�fVV�5��:Z����e)��m�F@w�N�G�f-nf3�h�F�,�~��N��mn�U+WN&^�v-$�o8*��y�S���8Z|����gMߗD�Fj��Iv�A60/uO��L!��u�{ID��?��f��h�P'X�h��-� #D%b�^3C�vx9
���r�a��o���CQ4��`7��L�:�7?��lf��2iM�(}`�a�2��( ��/�����$$*G�&8�Q	C�b�2���R���`j=�V���6��G�O���J&����Gx��永-h�r���J��8c)���Zv9w�c{`���]�Bca��}h{�����k�,be��ؾ����~.b���]3#���삱������׋��̹�#9�sǣ�;�e9�P7mR�-49�<�H!�,Ⱘ9!�û��s�iLq��}-��;0��j������?�6&�MD�D��4;�l�@m�k(Uۤ��d�A���9�Yu�F|> x��H�������<g��-+�p��BM����q�
�b/u뫢��$��)��w҉�Ij��j������]�m>��^�=��"?�`�J�\ם�܅�E�|_O~����XYqK�`���n��>���kB r��ن���_̲	�WSz?��PyX�m�
EpaH�ʓ#�.$��)��k�=$�B��ߖ���̷#r�w���C,��-�E�U�^D�$r#�N�MD�C1!��I���A�ʁ���C���;��5��:�	��Q�e��L��N�Ib��'@C��µ>�����q}����n���A�Tn�ĪZ��i	A�ч�P�5\�$��RB��kn�$��V}�;.a�*�*x�A�h�S�ÌڸjU7����P'�∏M��D�O|L�^������hkѸ'����N�E���M��厉�,�8��<�YO�-��f�m]�%�!��[&��VȱE��W����x���t����\�A�Υ�����]	�?XD�������t�~���Eb�-��
 �T���������m��Y�#����5s̤�#�*��,/k��:2�S7̳����h؊�YM������K#dp�7�*�~�!Ps��Չt�Ł�L˯2'L�G�Iz=� ��;�)�xQ��/�Š�¦V��ryjZu#}�qDT��� ���OFPZ����^/6�ڡq����ʨ��^�9*�܁ɤ�B�����x��#�/4�nKrNu�����=ʻ(` ��vs�^G �!d>M�:<�҇�������Q���d�����D���}���C E�D��e�4]��A�'V
nN:�n�\{���M'_A��C#�9��6�1�n��yr�ԧRw�Pd�.p�Ir���85W���x�>S��DIuz0Ґ
"�.r-�L��.ZK��L���ک��3��c��ׁd�UO�8��)s���N��JJ ���q��RW�f�V�3�e�9;jV�&~��,:HH���lޠQȅ	���S�����遙O����9�p~�A(��R�N��t��;�'��C"���r��ӽOwL�%<��;a,�����>�"���8�z]y�ȵ��q\0���j}3(��]đXzW#���\-���6)���*i���u�H���B�X���ʹ��C���tFP�d�A�
�+}��`��!5��7	����fV�-Q�OF��Y[v����3H�a.�-G��*i�D��څ2~�[.�ts�+��WĎ����	�>�`��Ÿ�T@&�6�x���;�_Q��cE.j�kx�WHZ� *`<ja^7'F[9^�c)	�� �٥`,��)�5I��_�pl.�6�L�l�+)����k��!�֮���[E&�����H�IWN��v�8�>Y��d�+�
%l�[���Y]��LN��M�a�-�ݧ��2�6�k�p�9���Ke8�f���ك��*��vL<!];A �@s��p�����cZfS#,M��g�����y����GT�`�?�p���<��>F���n½n���\��F����iݺg3_�\���\��j��	̜fn����y��N5�4O�̘�ʄ���z

Gcp�3�Ӑ�0�e^�,	��#ƚ��oH[��ƳKW����ŽN�J�1n���}|d[ȯj��B�E�cd�Ymmݺ���?��GN���i��<Z\^W�!��7I~����_8���4�T����8�q�Vm�/IX\a}E��1�LB_�
�q7���k�=�H`vZ@�9-����.�BL[5;"d{1��!��^����a&�\�ԹYh�-9#���5	�1��d�|�\1�;�e����x��A��p߼��C������/�gsl�C��f-JC}���B�M��rp7y�2��N4U縡���A��a���+5놜uwf:eI2���$SwS"�o���J.f�Q0d�}���l��Q<��5q�y�MW��ކ�mTD�ah�Q?A��8�������!V���}���4<�(�7h�Xſ���c���D�F��f���SD�Wg��Q���56`�rI��0/}�4����!:n��y[�l^�ځ�m�"��6H��t���\��'
iwS��}�T.i/֘��r#��)y"e���1��N}l$�6�����__�ӀG��_uFJ�v6������ʧZǦivh�<���O�.$�B�s�$��XQ��8H�j�%#��Έ�}p a��a��Ғ�Y��o�Pz9���x-o�}�!sѵŠ�s�ohS���	$�:���� M��O��[�� ����o�np(~���*�yI���5�� #&�s=�М��c6L�qS,���H}��R���O]���T��#���Μ��2���|ˤ�¥�cgӵC�k��!sDGc2+`&ԓUB#`�O-du�Uqjtc9{:4�M����]�H�I�-:C~�`E����3��ͼt�2�!���)�G��/����p�2WgH62��J"�3�$FFV�����q)H� gؚ�)�����i�U���4�
�Ù9��1/ܷ�L��;O�jd��������(��
4�T�U�Q����LH��n�.n����2�Ч�+~}�z�ض�,=�:q�����Ȕ=��Rɷ���v���z;�X��QIf�!s�Go!?���a&�3jfs{烦�u����Cz �|7�[A0�S�\��rFИ�z�i���)=���(�c��a(�QGA)J�=�G[$���0L��G�X�|��{B�F�
h����
�+}Q{}Iܣ�P�Q)�	���x?@��f�
LF�ʁ�^Z������JH5,��\�I�5��c��rq��hx����WT��>7Ļ�=�&G�~d��}4��EnL�:���W�Q_ψ����b�����k�vQ�O>���AN�`I��jbz��b���Е�U��l�%��o?�@~N�e#��A"�bOm+�Ɉ�z=_���a�F@���L��c�DS���q�;�*�g�T0�W�f���	#&B��ۓ8�k6��7oԡ�
[���+��N��D;Gq����208���)#Yp�z�x�S��[y�1uo4�u���lV�C���64�F����a��	���Z3��v�'Ɨ�/����j�x����ϊ���p �v�D�%<���4U�B5���+�z[�[�z�����K�C�*��[��)'�[�_�j4^��p����M�U u��͆Q	�'鵚8Cz	e�N��7���ZeeW���R7��Ȟ�ʝ���fZ>�Ԕ���$;�IQ˾���
M�0����I��EK������sp���`��g�j�Dԛ�����+}��9Ze K���Y=\h)(�SD��K��/��o���>����GCn����Q�W�8J��2��D�Y�@��,�i�	�O�V<zW��Ű�X�Og��^����|h�W�N�#�`����h��D暅w�������(�#�Z��K��2���8C�)6ߓ�]���2ML�y��(�o�F��;�T�$TЫ�,��g�y:$nΖ{>�q�I,	S�=�N�5;Z|5qd�b�U,x�0����w�m�,1�_��I����[tD�}k��c��?�=��-`�Z	N��ي��_�i�q.�����-ݶ%�����1�ঁ5�C�W
`�I�D��),ϐ�g� Ԃ�,ԌQ;nj?���2]��3֧n��ؒs
;�������H�`ԑr�/*!|e�"v�@�#c�;6텍��	tJ[mvޚ��}k�#��Te����8���x����ee%��'�2�"�U�t��F��1�1(M��8ϒ,�><��e�9	¯V�����!<Zc�����Ȳ�H�T�C� �Y��O<�⛑�Gs�=��k-W�6�pr��ڼ<Y�e�R�і��z���5r���
�R��(o�ڞ�n��M�{`�c�l(�����$L#�N/M^�%��8[�}���!��c�5S�<$PS��E�GE��D��kμ&O�Q �P?��whw��"��U_����ҵWC_���� �׀�=I8�յWB8]632���դY�3`�N�!B��:S���2`}I��m?��kx��ܩ�R5�e�{G���8� ���J^�ǧ�@����B`��^-k�F��SV�@�h����X��b����bJ��} �1x�Z8x�9C��-�xT�n�(��p�bL|�e��q�����=�ee��~�
�3�J�LMnH���N�N�?m�H�ގ%�GQ<�Q�����[�p]y�ƫ��P�����6$���{2`��U�����G#)�9z�l���,ƽP�f���"*�4R}2Ԁl7G�=�7[�,�C�������ͪ��$%>�����q��(�'��W�K'a��;��F�%V�������?H�JWAxu����Ko����} �y0&���H�i���qt�F��� ]79�u�*���	��*=EG�=�*[L��
|���uJ�$#���>�W[�ui�X,�Ŷ����|��X7��ĴW*=�N�ļɿuc컌��(����t�s�|mI��6�la�(�۝���o�}����W�&�R��3A}����;���	������G�ڀ7a����oB�,>�LХ"u��Q�~�����i詧�������5>�8��J���q�E<���"P�h�wj���o�M��ֲ��=��gkO�<��n���2��6��$:�u�s���A��t���P=�as����P�!>*��O1��2�`i��!]uA��,��p�V����(�H^�33��G���w`X;�f(��]^�:�
��WLV#}<
�V�w�6��U�'@��#ܸ�R�1�=ř����Ƒ�Lc��+K�kBF�`V���1vn^�Ǫ��	_����?��Th���aC�����t{-�s4ɀ�j_0g�<>u���4s�
?���#$�K޿��;���Ac��]Ғ���k,�$��qk�89�L�3`��4�\}����
�BiE�P��fU�*3���V,F�)��:/�R"`RTB���%�W��U9�Ʊ����[b�����[���*n��s<ώ6��c����yE�o�B�}]�I�x?F(�_B�!?qI�g��l2;�H�6�>\�	Ń?���eF�?o��:v��!�O�:����(0� ���I�p�r
� ��Z�J��H�7���q(�/��&-`��he��=��?�b���Yj~m�M?ݹ ��������>��3������)���M���H���9gAG���>[��
�l÷d4��� +h��1��3f�Y���6�a�'�5VCLb�P�S�U�?��˺*�1��t?�r��p:US,���W[�4��v'L�=�txvp���9�����y��4�j$Q����
|��.1.6�L.�y:��s�B{B�^�qY�Ĺ��
�:��%Uk°t�M�N
k���ϰ�u�wV���M�YC���S��aJi�[��j�H	�]�ᑱ�nsh�0ʂR2���8�$//�$R'�Y	���@4^��7�R����M2�7Bҿ�O�*Gh*�����v����!ߍ��Q�q-��ָSQ��o�����J2-�Ѥl��%�������|�Q@��_rL(nŚ��ӣ4qa�-/t���a��8�D�O$�5D�N��~��Ee���-��d��l(2�=ڼw� BL<��m����J�>�6����Fi�߶�ɪ=��<�I�dv�BV�0:�an��������U ��T�o	�# R��L�^ �~m]���"��`צ*�����1�#*1g�#������z�S�������8f��]>��~�� �]�g6����f��T��n��q2u�gR}ss��Ɉ�2�>�x�"�|��%y��^�Oƅ��L�S���:�'�V�H��R81��lqJS���?5I�����B$N�����	��~DL�\��g�l�rR�
3G�/\��(=�$�U��t)+���i0r-ݥk3R؊W#`Fպ<`%����[u�p�I���I�N1i���ZLp� 0�U'-�*}8ǿ S(��+���~Fk	�Y�2u
�QL�/a5�uh��#r�Y�Ú8�� j&J�~��i�_2��n�����ֶL�@�_����Vit�h�טS�}�l�s>ɘq�r@[2(��%���1i�KQԑv'�A�࿃�r�A�_�}IdCTѳ�$��)�BV�Z/I�?����|Rp@u�+�L ���".>�Ҍ�w�V �5,�Ƌ�ӂ�V�O�2g���7�:�� \�R_�)���F^�x~EP��q�Kr�C8��Є��v��O����x��22�m��5�.�DX�nJA�(����٥�d*�*�
az��
�����μ��sгMu���S�z�����8!�|� ����AU�.�J<a�� �Q`�{�dt��ţ8��&�]�xe�0�W�[���l�#[���W��\�hp���3��r����1��\�Z"��aܾ[>D��6$B��}��JjXH�1Њ3�J%M��r����>���u��pqI�����f�r��bD��Q��&OV���.l���� �c�JC��fF�Z����
;j�D���W��S�h^�!9☸�TMΧ%)�>�Y���s6z	q+�FT�]�@W#k7*����HÃ�H�9,�'���*}� �_��Iѯ9��vu	��YR�T��Q.'�5�#x~�x��Xs��0��4�%�o�`G ��Kj;ۃ᧍����l�Z�^��#�܅2^��"���+��=J,Y>�t����Ýc��n	.�>��SD9ě�fGQg&"���5�YeҼ>3��/�t�]�O�`��p&E���=��������'z��#vz���d�(R�{}w�í�=
�ŋT�p�W�*[�ķ�������np*�h߭�y�5�(���FX�1���#�_�h��,�%y?���m���<������ta�=%}^�Ĝ^'��ې��Z��l�1�9�d��*9�q�TSfq�ǆ:��A֍l6�5�%�АEB�l)�2�嚜�헎���zT�ڤ��ٷ�*3R���}����$��C���e�m5:���u�D~#�_g�K5�c��#A�h�TR���'6�3ޏ4�����<�(�5��#2�5��ǧ���_+�o=(�Ѹ6�g�ɩ�D0�_m�����p�U����F��lhG��li���]���F^���y�Ĝ���p�l��^����r��"$Mӱ<;!������;��f��yN��c��e���\Z���P�D�!b�ηO��}��KbE5Q��u�f�xֲ�G�t�Gk.�uq�9@&� ���ЏLt�M��zS�ΐ�� N��Δ+��1��R�. K��Z�]��iy�#˅
�®j�ϛ5ܦ^D�$K
��Iƶ�F�aڕ���s�X��b�@16���ʷsE��s<�=n��?oY����(�V�l?N�Tv�V��wUq ���2UT�F���s�����PS{�Q�*�i���6E��o���:��Z�ʶ�qB�T�m|�=U��9��/�*���{��KJV#1�l3�"�Ǔ_������
8�'�uLCm6��.5=b!W����-����^�!i��L�d�K0�}�k�#�H@��=c:R�*5���N}�XOI��d�-��^':��ڢ�|�
����<w��� J�1mx38��aqU3����[��ᤇ��|�����Ai����1�6�m}���`�O>,���Y�u�Y	��!��U�Xs�ZS/�Ѓ�r�ƻ��PR0u��<2��T�d+8`�a�!Ě|��ɉI�!�����Mu LIʻ��U�vP�7ׁ'dc�v��Kd ��u��-��1-n��Ez��Y��Z��A�P���$:�����{���-�d�����3�����ny/[�|�vطW�B�P��䥎5�������O���4(��9|�N���]���;���ҹ�,~4hz��{��q�%^��_k7����&(m�2護̕{�x�n٠� mGg�]V�|�7���_nl=�g�n��|�x�>X9T�ȝّ �)�Um�h��^{��P�q3�H��iH�����ja<� X=����^%�f&�]������Q#z̄�4*NiKXL��{�?��r��ݤ�CD����e���D>����q����GZ���)��uC.��a�
��2�����+�.����O�[u	Vx�`��%#l_��P�x�Ȃ8T�r~�J8�}��!;�h����%�Q@�̷V� ��}�'��K]]Igq�\�'0z`2��)׺�*�	n~����?t��8q���=�S��Kz�sK�b���������:���<�<'�,k��	?##��x��ѣ����X웝r|(ڍ\�/�urB@���������G[T"���.�gW��u��m]���%0W�V��Ę�B�`�ʠ��jzg��(zP~��i�tj���W%LZ���Z)�9��_�VGz��6+x���$�����c��H�]`hz�2��@�$�VTg�H�/�ߧ�_�qk��3�h�Q{�R����c��$uۢf(9V佅�Ƥ�����u|G��v	rp�\:H�l���Hq�ȍg|ެ@l־��;��P桗S���J�*ב~h|������R5icOx&aKq��*�_Ǿ�� +1=�+4�b�?������0Z���k3�d�bؿd�Y���rد������s�?g�ءr�� 3"�F�/��}μ}ț�V���Վ��pT	��4�e���Ȕ@r�Z�җP����E��e�ˀ������Dr4�Kk H��N|o��ĩP8kU`��d���w��1�w�����n�j��.ξ����Ӯ1.4�ſ��F���Pb~ߖ���@T�FQ�𠬷���$�m�M�z��O.*Mn=�I�\�����3a��A�DS��N;�?^tF[,�B\g��]q>b1��~d�
��A#�l�+�7$� �ʦ�N0T�4�y�(n���v[��7��>�lS��bݥ��0{x�Ŗ>6���Ù/�*ze�I�E(ʴm6H�G�O'h\������Al&ZRܭ�e�KGY8���֥�3��a!�e���^\���SPt|�[׵��E廳Ͳ����l��.Ҿ����)��	�5S�j������g�t؝����($�8�?΂Y��tCk�!�(� A�C��e4|g $��b6�����y�_�mʱ$(�jN�E�b��A�v\uy}g��0���8���@bԘ�tu|6B���ٷ�6� 1躝�](��\"u�}���
��z'����=n ���/��z:QxE�e�:��=�+�l���sa���c�I^vi��|p�ͅGl���H��A.�G+cb�*���y^~�f;I�ȽJ�i�]<�<�.[ �q1��u(��EB?���E�U��C��RڕP9�lJ����X��-mE���F��V
L\t��]�2�2�5k)�X�OB
h�×'�2�����+�e3oDd����n�kdO4,��}�3���r±���0��m6��o[�*_6�N����#'8<�X�3�l���y"l�.1��#R�g���9Gg���f���؀'�⬢R�)�߇�FP�i��nظ83#�J��f��7kye��Ҏ%!�-��b ��ϟ�ݤ1����1�4=�l)h��HܭyVZ�/+G�&�:�g.$@]Ʊ�*9.GC��A���C�����"�;)�}Zq�C���1�g|�P ��]�u0����!t}h�*�v��uT�A~;�:\�@��Ӣ��Mz�v�p��i#����U��)#�P�&d�E�m=��t��e�U��
A(�lK��sfo�`�̡���:��������mm���EL�
���x.��%ܒ���'
�7���al9M�!����9��iĨ�E��9�XP�z\J�^���R�i�@g�C��s�������'���7���C^ZP���ur ~L��BC-,�[#z�?�1�L�':�L;��)����R�S1�4�ͺ��#����I��N0Wg�~��v�5�-bgL�_�`#�C�֜RO��{�Ҍhi������ܱ�v_�~�����ؙ'�AE���'M~��t��\��]��T1��y倕�o�D�����NV`#�zG]�-X#t9̈�>7pnl
��r���m��V��a�X�U}�G8�p�2�p^�U�ӊ=��U(�(������t[��f�s��n���-�[w�?��1ט���P,���ַșyΨ�Z���,�Lbg��8�0cz��B͊ӱ �86o������/��Bի��u��?�[�.A֠-���,�7	j�?�u�y7�
�t�/�s������;Jع����ӳ�(Ȍ6)�������=8�����0{� 	�����b���,];�קa��$���m��S��<½
a$�+�<�KV���d�r�vu�(�X�_7#C!�ӆW �^�+���ؾ�d5���<� 
����I�c���^-0m&��[��̧��`�3���	�sܶ�	�~V�����nc����ÇU��ެ����ox�)�W*�����p\�5��.Y*�ط��ʻ�� �2h{�J�d���6���TXg�-���Բ�VE�p��0�c�1��hY>%>`��i�C^g<&����d�'�Ra^UW8�=wԌ�/�>%Q�_rQ�У>�_������������ӫ���~e�w��������x����B����"��:��JT_��a���t�Gl�q�4p��a'T�5��S��*�J���d3�%��u�� �T�i("槝a�hM@_���+�����l�Z<_�?#w�T��o�4X?��&?���@�	�XkV�~h�õU�  Ջ��\��u|�c*D %,��=6s?{��o����a���9Ց��a�Z���	Y.�i�"L?nB��@�\Y���>~Q.�)��Y<�HM���=i�)���Bm����̋�mW�	��Y����J�K0�)�	�ő�����8!q���s-dR����/�*�E9^��j]wc�Ϡ��O5TNv� !#�SNJQ�^�!:�']7o���}=[N-9�RK~ϣ�d�Òm_��@T�0�	{t��W�Ƶ�BLM��F^g�Y"��y+�����|}��ա�r�G�TR� ����61��(��ޱ``���W\!�d�+��_�"�+�6�,���	G`��v�%#����$7�l;P��}�,ػ�l�s�z�
��J��C�%���0cZ7<qQX|��#�K �R�EOԗP,��f�k~������ʃ��xLc�\�c|�Ga�-�aP$�Z�1]�K;� j�]-~������w��!���.�O����5|c^E�ֹ[�M�أ*�NX���m�;��-�o8��P�)��.#ș޲����w�c��;��Bl�����K�ݗ_��o������4�I<�=]�"�B&�sx�}R;"h�}�w_�I4/�L���B�t	�J��ge����
Xj�+ns���}S��mB�{���lwf�� |����4�f3�-:�T#���������p�a:3�Z�I�� `���G��jsǹ@�Io�x�*:�ww���o+��b���TT����E�N�����6��T�G`!"�#B3N�nH|��C��ݵ���W>��+2mZ�]�赺�W�
�uf��CF�'ޫ��3�}4��������HT��jWB�����m1��q>Y"㋵H�9ގ���]�棳��v��	�o�T��E=H_C�lX� kaRA|�e:��n�� >M��ā�%��u��m�U��9ia_��K�%��7�硨Fo�X�:�]A{��5�K��2>�?;	QJ��)xs��ݳ�pH]d�1TCY��,D[�� Ipc�t�5h���/�h�����a��y��œ�%,��"�'-z�Ȳ0X��3��, }*�ԛev�u	g�Fn�䃿%���?�&����ǡ��Du�^<��͊��m�P'L"�aK�����udb�J��D�����,��0i�����X\�8��v�?�Ɲ�MB�8zIB���n(v���NgJ� ��F�i����>	����YCm{�/��D����rs�;�O:m���3͌��%�*?�O�����e�lɤ���ظܧ��ą)�].��MK��Ѡ�~M\���4R)ʕɵUi7ӡ�`��9��iL+`����(x>��d�u�f��N_��.�b݋�(+:R8��7������������M���sŞ�
ؙ����7�i@& �!4�+���5��P@��T��_oJj��4��Z,ZAt|of���n>ˌ��R��t4J���4���"����|鵫�_������L�c��l`qb�d��43�f�3p�Cs��&���T>��řP���?C���O��U��0�H�J�}uF��泥�=v����޲�W��eQd�rA �
Q�DW���5^�Z�vE�զD��2�mT�I
�d��i@,�4�d�S�;=�p.�9F['�c!�޽� �t����}�"��S==�ڛ�'�U��Ϣ0S4i�� >�Lp?�W�J����@�Ք.��2+��`��nC��a�X��܇Qɺ~1��,+ <�ϩ�����pJ��7�=C��S(��BC��重��%�춹}5�;��`���qEWT��N#)��B�������`5�`i��Q�ݱj���,8�!s@L�w����t	�����
�+�V�=Y��U]sc�`1�?�k�����f�Ԯ2�胏I}�w�;|��"���jί</���,���p
"2AB@E$�,�ű�b����v�l�/L��ꑹ?R4,����v�XQ[fP1Z���p�m�ᇭ�;X�����}>"Z��dl���V�@-_D�R�����)��xV���[���f��Fj,�Y3�[�8�@���>*�㙈��zO $*�}�� =@7��1S� >�zҩ�N�ܣ8���|YH�eO��_G-��R������D2ڮ�n.��ɢi�߲D�k�c0��]Ja/B�|�j����+U�}#�,n�("l�������\���
�i�Pn�
��"(�	�KRH�����W��r�Щa}}�&8��?x�U�4I�Z��	�{�y�k+����f���D����8���[�oB"E]�O����}��0��{Ս���i�k|p�7tR�䎱I;o��N�bR��:��@xU���'���'��W��:l�	�Q���<�v�-��#����,;��@�#@.������@2)L1��1��i�m�����0C������9�99�e�LYN�(�~��f���$C<���?�b(�<��53�;�Qh��j����#vH�(;"��+�u�\���H�q����e+da�EF�0P��7����{a����(���~��z9K�%��]U�7�cf�]�7�fk=�aH�aD�o#�����
n� 3����oMHh�H�r�.J�>��8���DO��L��O���g��ۻ��3k&"٭���s�gA.lޘ�.�T�A^�-w]�4B��T�:.码�ݍ��x�m��!�E���̵Q���	��e�X"�.8�Cm��٫
���%�<N1���E�PJuk�V��N#.,�P�q?����V]:�3޸����Ta;�����Y�nU��eC��E�
Yf�g�2�q���t3 Zc�R�A�Lm���#� n��������HKZ�ɲ���Κ�&v�T`닇���=Ν�� 8��A��Y-)��������h�_��Mw@c�D��~_`_�g�_�,�a��"����f����9�&Se��뇄�VR�ߏ�r�ZN���v}��� ��j]�=b����`�WZK-ԒiĶ:D��/�P�G�Ѭ�����H��Ԫ9�$��qx�
Ēw,���9ܧ��wD� > ��t���d�`��] �|p-[k���� �c��g+���4�/��"�]��
"-����<�q�H�c����N����/HV;5�B0u��B���^XF��o5��R��+Y�.�pT�#���ϧ2�y-�$�(
��Z $���N��$l��-�*Ԫ�I�����2I��c�@
��>�x@�
Q�7֎n]�Y IL���8A��'M�ՠ��L('���ә����J-E=�_@���4��GA�%z�ދ4�;�4�&���) "M�ԓíQյ�}CĮ��1�2Ɏ���3�1؉p������z�U�䡩 EH5�[������� H��#W����2�O��-E�����y�86�k�#0�$e�f:0x�n��5�ȯ�n��c�����m-�&���N�!g�w
��\jV�Q��K�8a8�3:���.H�(>V䧃��?��D�Z��n%�O�)wLCU\.*{�+��	sj��p+����j9��ϭ��8_^��t�r���Y�;���0��xS�-DS5h��2Y�::lThS?&��u��3� =�.�
	9_	]qT�S�,�&���:��BDN�ָ�m4��D:_������![|�Q�""Y_;d�E���XX���2޽@�|`����U|�����eթ��`-4�d{��y��̹�+|��!�
�б����4f�Cr���-�����c�����:5Y�z�:�8@c���hÖuδ&<�#�Q�(�Q�U
���Kј6I&D67V6Ϲ��"b�cy�#O�n��`.%K�щl�	T(� (�N��e?��-�4I6d=�ӕڀSs���tY�Doь!�*�\ǋX�v�]�}�#9p�����&�,DѰ��B �5�5�A/��6DTNg?� : &�@�͛[aKpaRn�Ŷ:蘑mF�����:�������/Ǫ�%ou�X��?E"�a�P�����>�VN�|us��w�_-x�ҾHg�I��I�]��r�� �nO@�-\�Fϒ����a�$}p-��X���Z!w�C�du.?���  �|����k����R�ŕmu1��^�Anۜ�j�k�x��g�Lk���������ya3#��eJ5f��o'�\h7�b'5x4�ș�ةKɛpo�¥Ka�Dڴ�4_^��%���:/-�I��}_SX�8ǁF��Q��g��x���a��@l��f��kpz�ж��[�?��sqᛊ쥷��b6��r��D�d��5G��F"�E��^�Jzw�]�~��j���#~JD�׳v`�*G�J0J.����D����5"�k�>�0��N��[j�3�8\���acN��6C�.���j���qq|�t+-/K=	�d{���G5��77Rb��v�'���yw�^�O�h�,��0��g�'9�p��q�mX���`�N�o�O�g�*�*���!N��L�쪷���
�w,�?��r��i�G�};��(7�˟�#���^��Jy_�C����)��m0�����DK��12����+� �5Q��=j�Cz>�n16zQ�!S-A{�
����Uv��[�_S�*3}��=�
��+�`m�	}0>2� ����J�D��Y7���;ǇuZ�ɶ����w��� ����~��*t���Н#�彧��ހ�O��~�[�p�IU�+s�,�X��r%��ܓ�Bd#�X�Gr����q=��:��b��y/�rU+��Ƃ!���0���3`�# ��� f�'�}��Pn�;x��c`K�ƥb����C�� 'i����S��o�SC�V,*���}.���en��׈�]��y+OՇ����Gj�rF�/�Pj�sy�k}pp��Lxv۱Qc˞�������#Oc+���!�Vl�:�m,�eBdXN�"d��Vu��K�\s��Py=V�S�M�)�Z3ܿ�Q�}Tʵ�ow�	�,���#֞$ �ߝ,��\�A?�j��FN6战��Ս�y:vQPG���	�B�՚Q�=�乀��7�]���ޢ�M���/4`>�f���	��{�I厑*��?#��Q���&�}
~}T�^E{ki�eBjL�֟��3���9��@���O�9^u{��;e���Ȳ~,�p�Ή���X憢�P�q����J菔d���SF��@���f�(^�0Yw�F.=u������/�׿����#�Y��}I�\8���b=u��Z�C�"ԛ�"��N2�<<� |ύ`ѿ��&�	�]"�ܐ��F�BV�	c��h �z���ʿ)��.�O#X��g6�D�٪��Z^)@li��қ���vfG	��i��3��y�t����S�Ƽ1�j��~o�A��#M/���δȂS�<#����|r�׊�����P9���d����ѫ�wI���ν�� �Et-\V�SW>�"&�<�������?�Zy��`8��>u�h�D`��hK����>�� �␧��Q��G�Ʒ��Z�&B3O��]�������'�.�/��
}�I�y^��."���(a�/w�Bwc�"g���E{5�0oƺ�f3^`��2D�\�E����q7:k&�^��B��E�͓/�,�`�ѹf�΢6���wpo��7�2�l�B���pY_�Ҫ���0;~O��!F��K�͖�����k�kxn��|]���?�e���)�L�@�����b�ð�o�MD�yL
�m��?��L�SD�m@h��*�͵�)A�{p���J��Mr�/�j���U�X�M��Yk��&m����C�ᯃĥ��*.ʋ��K�Mr���x�;6��O�y>�@m�H��&B��W�G�+��>h}�;���\*c֭��%��x�B��r	rʆ��mc|�Y�t��͆�ư�Y��|��9uu����ث��D p��<�CIx	]�3��"Vq1�o���!�٩����{�h��GU��#��5��qj�T�f~y�0|`����	#���ƥ��BR1���S���1;�l��%���eL�67֘���1j�S9���<�cn�T;�j>�pF��^����Ĭ_2�B�_9�|�4������Hg�I*V���I�P��Y�򝔸8���^3�,��ws�w)?_��b>8�����[��tn�o��>C�|J����2��T���&��y���Q!��ږ�$:�o.����9��!�W]yv�����NS�:Ť�]�氃!��j�v��H����b��j���9�� P[;4���)�m,�D���ؿJ��;p��F]/��4�����f�@E�y�b!P]����������^ؼ�����H(ļj�m�l7�"�֍;!�(�М�W����#��|@�u��u��jY�l|������WI�7��z?���c'd��nNk�R��4��ұ������i���ZkL&�&D'���G��_tLN��&�,icc������5�!��Q���*�\W?���������iO|�X#eM��|#�Y%|�����UÖP�����)8�'_^:���e}����D8�n�}����sc�-=�4hf���mn+,?#�(^+�S�Rn��*��"?r�::�n����a��6rx)-��Q�y6�� ��-�sgJ�����a|�zRdG�&�H�1�زH
�.P��+�;+͐z2����ᗐ�`\%�fƄ�����Z�.Ґv���(�8�p�^}��S߸I�&�?���c���9�V�t���w:��M�����磓�u�  �{<*��/�(I�H�����"�>���l�>'���뇿~�����w��� u��'G�r��\�z�� )m�ֱ�2�T�>�{����%Qu�qܪ蘇t1��]@�4��	ݑ ��Ϙ��G6>%\qQ6[�L7�<х�����Im�1�����ۮE������ CΘo��X�b�xrf��9or[[��&�����m��/�B����-Asa��C+V$�&�Ow�G�^���K�E�)V��z���H�I�b~��*P�k��taB��綝�)�""�0q��m9�a"��7Fc�#tm{�Gb6W�6�|��6�SGU~z	68\���6��ǈ��wH2ݩü_�:��)UHkᶜϔ��$b�F��uvx���j.PݞL#�������7U�6#u��N���23���_��) ���;׉80n|��=�"(����c~v��A�gZ�V��~���f~O�GRS�ى�����sgw�MC�߲#��Nr'i��,#�֤���2v�5�˭$b����6��f��4�B�� H�(�aq9�v �8Ҭ5\r���Z��:~��@~���"�Y��3��akFO�} �����|����x@��;���uHǔҔ�TY���#
}�q�R�������Q� �wI:�t�������ÿ��9���^(��ؤ��������ܜ#t8���I�E_~�������ܱb�����!|��U�GS&0AS{��61{@���9����_j�?�!�.�*�]e��)�`�vQ����H䥵�]�;��Dx��]�B�+�f��#g���\���]��].�"F�H>�]1�B'@7^�^'���'[Y*X�lڕ�D]���N�ȹ\&��Tc��>\&I�;P!>�M� ��g��u��-(�Kw�H �e��n4Y_�AI�[���$K=�~P��ؠ8i�fRܒ(�ܼ�4枩�o�v�F谾~b��~��9;��0�_��hp�jt�
��`�� c��
oa���D9W!���B�r��π�u������պ�4Z�;��I�$��ۻ�J#���v7�\��k`��+@-O$�[�f�ObB�C޹?%%��u�<E:V���m�M�8T^o�A��2tWU/p�6Vُ�n�[L|Q�XCq��B��A�D�2]�����B�'����OD��QF3�qѭ��Xhܦ�|���#Y�0`��'���[�*����k�e�oh�Q�|i�t?���P�|�nu�RV��r�w<F��q?�`�`�}W�"��*(d�w�����~�Ş�!b�F���!>���0/��'�Q���F��7�J�?z}h���Y������&��_���!p8�g�V�np�o/��mFWwQ��8�@><�#���fa�_��O�a��qsUgQa�ܚ�m9� 6���<������a�s�y�j�ZF�!uU����^hb��n�(���]�X����wl�Af/��2cp��C��c*:�/1>�q	�b,�ݶ�)��@@�!�Ns#�o�]i7\�@����.B�jӸA<��A����y� �@��gv+jt���Hc3>����Q���h}�&�L�}ô{�ذ�ݷ�6��!����E������5�fu�Z�� ��tdew9�������U�?�PL������;�F��qU0Y��-��T2�fhiǌ��d������[���^ϊ�õ
Ɓʀi������l)�~�d3ݢ��#���հ^��|�rqv��y�;��i`GQ�D�u���$�8��vq���4`�Z���N~=�:�l��*�q���Ƈ�/���M��)���vd�����c��l%�� �����'�j ���NQtU#w�k����X�H�-!�»���ea��H�]e�� 5c�������C�qyX}	�9dA/�G�?����/?O	N�����*I�^�۠�L��)���y�}'�'�r��!*�v��)��k&{�$�3-�[�̄���-�h�ܨ�Y���6AӌO!�o=a�8���e���7}W)�^�<d�9G�b�e���&�+\o`���ϴ�9�_e���'�̸�d��`�1Ʈ�~�Z>i�=�եyB��m:k|��m"f�=S���=���r��`&�<*�	�I~��&���ܩ�A�e�%����
�<����^���+9�*ޝ���x���mk\ٯ��f����N�c���ne&>�R�{�X���%],rGά��	Yw������T�1.;��П{�-Iz۠.�*�L֥���ɧ9Nf�ǁ�[S����'�O2y�k-4MD�o���$V^���9^խ�LHHI]z���{�����[�ͧ?��#�9!<��B���A�$�T���)�L�A�Ka�b��A��@#/5�է����S>o`��v:�W������L�ep�Ǜ��M�������Z��74FH��.fM������Rƛp�]���лw��
�a��,�W�Ϳ���<˛Ln8v?B4ׁZg58+9.ێ|�:G&ߣ�Ȅ��I6[FP�l_x�7SA�羆�N8��,׼1H�������W�J��F��i��.U��
��׉����U5��Y�S)?��j͘��wڂo�o��j!e&��wW}��^��y�$
hfTݾ9�/'�Lbf��W��h�h�Wf\�7i�gX��#L�ꕄ)�vB��&�{�.|�g,�w�����$�'���k[�A�L~�u�'ޡ�.�������"x��l?!��սRT-��]i�N��`���4�̮B^�E]���A�����]B�����tFP���ѪO�DFiE��@��Ӳ\.�\�֟�yk�O��_��R/ ��Lp�Kbr	^|���R�z�	{�X��>K:� 5`������q>:ݔj؅"<J�����IG'��M�ab��H�]`�����2?+ܩ��?+�8p҇1 ~�Q\d�^��yA��M���k��M)�@��MH�.�z�C�}m�&�	�ߵZ\ƻ��X��P�gk�/:!t��2��y��`)�6{E0����Xz8���X4��L��[���f�h?A\q7��z$c��Ժ0y8�#<���ʲՋ962��*�
�	c�>��HLvt��������A�¨�?[�#�Uj��Qen�R���Bf���b?2��������s��
Z.�
�h��ھ�K��S%��OC��x�?\S8��[�vM� ��樲>�Ó-�l����%�-���ɜOH]�v�}�q|�.�/PD�[�iвy�'��%��R��]�ʚ�X��P��̱!b�@:G��~	3��ϼ�J�	���0�4p&A��y��܌�z���A�C0�M>�hN�x*~� �Q'�(�Ξg⚦�`)H�pЭGԙG2�$iᣐ �a}���!��NbJW?�.>�.6���G]sP�U��r�`��4�:�2�n�ך���~�qɩ��6q)�h�j�e�Ho�i��V79SR��.����#����.˧��$�,��l�����!|������!Z�W�魃��SG~����}����LI>�ֱ��C���B�;�Hb�T!�Oq��_����CQp�?V�1��ۦ�r�5hd�̔��k!��~c�يg��ɽ�|N�t�\�a��T��tgͶu�w�6*�t:���%a�9L�s��JzG���	P{r�\�r_[@�����iP��Kr� ���p�	�Jɥ�����0��
'�:�b���#H�e�"�Ԭ��;r_�t�d��3
�R����S�9'8H67��Ȉ=ް ͅ4���W�끈�����.��j�<�E��wvY��ռ��1����$��,��l�G�qR��;)A]����⣣b�]�H5��'�R/u�eRz�J�L�A������=�5Wʋ͗��،���F����o��� ����jo�g��Ɠ��%u�_v�mc�T�����˻� �����qs{�Gg�;n��Pd�v6�W��07��.`LY�a1L�&x�{��Rd��$��Է �g�璾�x���n���[����;�.}y���p��xс؟R�pJ|l�S��CLO���kي��{��h�.�x❢1��|���P�4�98�M�d�}5G&{��kL����A8�-�� ��P	&AW����0��Q�#})u�g�{ކ��[7����_9��\x�ʔC�H�%coA
�6����Cz�L!�������,d=��S��>nyƖ���l,�玴�-�YɄ��)�aF1O�?Қ\�9L&�W^��AO3�?��p�t��
�ч���D�w�p.�kq�cd����M��?��͉��dQJ�2H�v��r�tr��1ik@42���Y���/Xkv�g��PZfk��Щ�כ�ꐎհ.���]F�0���Q`�:����w�"z;nn�j��`��(�@0��w���7t�ő�)W���y���͔H\\��P,Ý\̳�r-�ᕂwB��4'�� F��8��Y!-��L��v$�B��x���^�v�B/�*��ぼ)� �gb�#]�0Z���*XfSj"/x���g����D~NY��Q���8���C�4�V�y6E� d8w�JV�l��X�c|8Эr>��gJs�5��:��w�#�5��m��3|Z�x�^W����~ :>,<��{{�Ș�>Y/D*M���M��o� }KK Ѽ~!.�x�[��%��l�sPd�إ�b�E�,���/m`t\Q���߫)0���^�z�Y��;�a��6���RD���cq�{(�X\���5���s#')��7��J�����?5�6W;9��T�v��0��!�Gh������%�r7|̛�p|�ChcL�5��N�圼&�"B�Ms4�����NB�fȓK�5aP��>�op�y����u���%��?�7cڶh�,yxd���w��?m�<�M�ūO]3�D�9Æ���˟�����v�c	h��O�y�K�����Is��6���*(��Q���$4����oEg4bS��)W�m/��+��懪��¬�9��9�m��E���d�;�3�</�Njs�A�������6|�SZh}�RS��o�17o�̤�z���ju�gqL����ѱd��f�eA�B��O�
���jqIGl�b��⧊�)����Mqf>�GU[��t�8�`��zJ��?���-;C���J����ɼiD��5�uT>B�ê � ��e ל�Q���ȧ�%�3�\�X7'�sM>Q����� �����k����2���5��ؘ�6l[�����["�	)�e���i1�N�� כnx�XO��Y/v荅��C�9�-���$_9�N#l��G�90��J�[�	[m�U�tqMJ��I�� �m'b��S?'P��1����W9I��{G6S�ڇ��]�j�1��`?MdZbZ��m��y{����S!q%�k[XqU�Ru��z�̵tZ�ˍ sm)H��P�6{�k2�hH��OZ��x͡Q�	�j�l�F���0���,S���9���9+Q�:�3���Lvj��8��+A9�C��\.u�4z� K������G9yw(#���v��! ��wO�Su�[�Q_Y��Z�Y�x���-`�_BX�eɲ}�e��ZP�Bb|��f+N.��9�׻�}%�}I���A����$O���7� 2��7.�9��L{ß�%f��&Uh�ff���t�@���8�N���vQ��lG}�tO��&D�ð�T%�W��dtZ�(���B��͚W���+v��!S"��Vk3fՔ��귿5��p>����5v]��Å�l�ͫ��s�L��\J������ξu��>U;����*+c��BC�ى��p�U�B�t\�5���;��6��l�eM9��`�I���YjNN��R��f1[��X`3['�f�J8���l��#|>���k&�u�ޱȊN��A���1��gf2ȑ_�~�o�]����̥WK4߱�`l�4�u�����V�j��W����=΁��N�ډ���m�
�� ���Uy�N�V��w�ۉU�
��S�"��vn�+�(�ל�� /OݖZ,�P|"���Aƺs�xrbH�A8�Pa
���F>���Ġa-@&J#�.�;�S	�Y��wû~6���X��W����s ��h�8����K�Fw˕��Bp�a:����0�.o��H��N��}�dd�J菵��53�C���L.�k�k+���e�u��&��13o6 �#eL��,&0ƤK�6��$4�P����	s]x�}\f�;�l�JUxl%���K������R���3"K���yp�\Ś,9Q�,/�yܣ�T8���Y���Q�=[A�=b�Y����vk1����}�j��'�3Z2��3O�DҾ�l��F NorF �vY�i-�b����nx��y����
�C�]3 ^�<@�4k���?YBوY�,��i�T�d�C�Y��	P���	�Y�Ԁ��
����
pa��GF�
(VP��XC񪍓4�����SE�}�l{Q6���Q����'`�H�˧��ri�$�#:������Y��ă
�"���|�O��u^��D���׼F���L��f�4��TĜ�S��LR��N�)�0�|9�X!�� ���C�O|�!��Nu��H�:kr7LI�q��U�q��af��V"p�7D��\���z� ��C_��1	J�{�Vm?X�����&� �!Խ����Ǖ�, aX��?Z�s�D?y,�^�8@~	���'�ma�����[U�H�s���c�8��P�:��a\2�Bo��8��|GTt>���`V�-��4��R��ᰢ!S�D�hA^�+�r�ӡ��Ǜ�)���e�WZ#��!M�(_Jr����6E{�7��t��~C���l>ȗ��A����hE㕻�?ٕ��4���.~��O�Y�U�Ԯ�3G;ж9Np�e���)�a�J���u*m��+�؅p�W���X�s����P�FCrW-1�RVƺ����~����������Ɖ!�	��o�=�����v1;꺌�J�TB�~�R�3\R%��RŠG)D��*@�ɦ�Ŀ�x��G �([�vV��f��{�@D�0�%�����SId@�_s��	;�i��t�C�ĳݎ�V&�\!�FV�(��r���P4�H��y���5&��;�N�o���t�ʅ����G.��(����'x$~����BҔ�P��]�?�nF��ث���/��N�[#��B���Q���[b���R��v���xǚ��z�ߛ�s�f���È��!=Q6G#�C�}.'ɀ�G���Q�8����"̭���+4��l"�n㈺l�
~}�1n�ޛ������L)tMFj���~?5f������eq��G�T@����Y	�e�#�M�`�����C�1�ɷ�byN9�8b�8�V��'p�WU@��1�GL��� $�����,]5bdі'i]W��`�x�g�jJ_�'�:5aaL��
��Mŭ��N^yNiEw-�ĭ��RDwg��]؎NG�s��M�$�8h��x���}�G��ӯ�N.c�"QN׾]șWe�$��ys�~�FÃX�������}��@�k=*9��H��i��ghT���1�?��Y5Ա�($�$/�PA��O2S�9���%��F���^�#'+�߻�M��j��R�������@2.`�o�Y쮙�C���(o�ĺWhU�|��@E����<��V~�*�ǹ�6�.E+O<i�u�6(R(�NpL� &�d��o�[]�z�W6W2���Zk!���qY��?�/�xL�7���%�P^ˬ�yw�}l�B���}���xgk%N�*o�M0jkK10�/� z���e½�(�T�OR���4Âx������!4�� �	:���u�d)9T�+�>J�f�����rvR${|h��"-���[��ɚ�����t�r�66��[�	�����!�A����<���UU8OK���z�c^���v��eܵ��43������������:5��`���q|����7��-:�����ɇ.23։cHh���>=������R�b�Ĉ2C�2w.�ju��7ֳ���/`i�=q��QPt�'`�Wv\��,$���dZѢ�r':�M'`�٫c�;�S�L@jgy�F�EA�Ne�j2�Ol��	>(��`�6:�A[קd�U���H\D���{���XtomWgfyO8�B)u����;ۓ��H#� 2���z7�����b�l���RO1�����ʈ�J�BI�OE:��[{�����|<�U9��ŷ��U���PhnDՇ;e�U�1q���+颊�3��O�Ʊj-r`.#���`9$�@��~7��cM����K��9�E01���I�[I�ƹā�U��DeW����͓->)��[7���I���@�1��'�x��ژL�'K�1zۜ�qI�r3��}8S�  `F�`\���R���GV���1O�p/-k�R����X���۳�Q=�V�/��9l�V�EO��Se�Y��'9�\Q�~��K&T�Ž\��z&���|��Ƶ��t}f��ᯓ��!yBN`���y>uvv�*Vj�A��Lf.��_ŪbBO8ûf�}��8r��웉1�Nt�Q&�<����$Gf��ώ}�۟���ߝ��w PN�o��tg/��1����֊��[�1����"@�F�*�����U��J�����>pG��j]����M��	.6�u�l�-9{u9`M�&o��NT�pa�6N9�֟(���kl���?��rf���/��(�Z��T�b��zD�̩�"��;�=x��Ӡ%�����z��,� >Z�=(�W��c	�}�P��qa$	$���G�qom�NڗX�~8�ˉG\a�@,�*ί4o��HDngN��w�+�Ny��+�|���ÿ��Q\��-�̝�rm�49U�dD*��D�}vs.�ʷLM���# i6��p�6�["��x�����f{kY6�������:��-<p�$1��1��������	UU��E?Z9��Lto&&g��$�Q�Sx���hO?�������M��bw;W0;
,'��?��8=�+�X�8�!cj�7<���s��ܺ3=M�R�ߥ�c����vo�l[N�29.����<�%;��@�K��?ф�$_�xC5	;����g�&���Q��h`4�����&!V��i�V�ٚDZK�'%Y�κly؄ô���Í�]�2M�_6� ��p����x�P�֑����H"�e_MZ^^�GJ���~ÜVj+&�*�9Ҭ�"�T��}</D�������F�U#X�C�\�~�E�.t'A���`�ywz����4 �r1ؑ��@�ؼA�uJE5/Y�_z1�a��T:���t�jђ�����U���$́�,ɞД����M��Z�dñl�@S��T���UՇGݿ,�ۇ�&�����	D��Q�(��Rf�b%Q4��D8gM���t�T����w�?HQ�{�1zkF�����R��A�%�Ut���ޖ���F�"�+�(�5%���ƠT�n�~��������һ��;Vݷ��6�f�$��.�l��@���*q�� 5%
2?D=/����I�U�E��G�Vj�6&[<�=�<�:}輊f$k攠'����a���m��� �p��:(Ӻ'�C�A� 1����)�ښ=$Z�B�\P��<�NR󳫫�F�e��.7{@�A�z8(f5�mɶ�7����2<�v���GbY9Jm�"�}�\������	i��N�Ag�����&c�f��������DM�<�hK�{�΀"VD8�����յ���B�46[� �Ԃ��5��m�ܓzA��'4R�Ӻ#���pS�Pp!��4Ѡ%�������!��o�g73��{���Ppu�и0Ћ�P�R�1U��6�ƣ��=���ȑd���nkN� e��h�:= Ȟ���^O+�>��;�!����7]�(fF�2c$l��i3[���W�oT�.�����H�Zywdӂ�#�0�1e~bH.�'�0 �P�"���-�V��T��բ�Qo���!8����1� f�[#��D=�d2=UO ����A[�>�'��}OV��8[�ޢ����-����`������QH���@X��/�g���!�������4�'J��m���>��aNpZ4h7�p1%�U5|��Y��^�S��ɫ���w-�eB>�'���~�C-��m2���y"��2%���3�����%;yG1 d}�H�T&��xbUB�T�\� ���Y�W}�VyE�&}�Hy��vp��DI�����@���jm���&�y��3@h�;���9"���lJx!c�9E��]X鬋���E�}/�w�^��gj�J��i��E���vb���RK5'��)��9R�ʂ-�]�|<��n�Q����+���ͽ�1����N��N�SR�`1���E����m��o���'���0�^(�~::r\���-ȓ��+��W�_�]��T�y�)fq��JS��B�(<�?l?A@�/tJƺ�ԗ��	�=0|\l��!}��E̚���3_W��(ӿ��"���Y���10�l
ti� �ҔkxA7:u���~8��1�g��L,'���H���!��N
Y���ij��{���~�Ǎ�V&���Pc�����_���:���=�G1FT3�BHr٥�g̬����x�QB^Q%/�R�@���8����?��H�4���T���S$گ�D9yL0���gKk�t����BW����ʭ�������_D6�W��BQS#�]�qG��\���L1���i�5����yW#�v@�>$\�)��S^���m�(&���|�����m����ʧ��o��OvewH�i������iu�3:�;�k-1p��"�w������w�_8b���k�'��ݮl�E�����̪,/�[�fGR�V�rW���C�P�c1a0e��	E�N�$�R��@C,�M��!m���o�L�e�>��iЁC�]�+�:^G�8`�D(V*�_q�w�	��������m���E���R)��a������M��.����U�?�?��ِ�%�o������G��;ۿ�^�R>Z���m^�IӼo��� ���3*v එ�o�*���)��`o��*�3�F�\��L�t��Z.x��jBh7�]M��ԵL�O�h-��Ir�g�E��X�4�C ��u.�h��Y��S�,��.��wV�y�F��A�ЦϠ :�'�Jw����[�l�]x��(S&��Z��P��9��/�"�PQc6:��tZ[�7� y�R��7�h.:@���a�?�[��R��-�]"�>�fX��P=�Z�������<`HsF+p��Ԝ� dt�����VB��i�}�S[�ã��#�?����P��T�`��F�DF�q�ר2.Ln	rB{TW���c��Ȁ(���c�����82�"��سȺ�r�$K����W��SX��΃����E��h�	'�Im��y{{�Q�� ��b~T�!�;ؕt+�%���Y���Gw�Gߪ�ڴm6������0q�l��#�x�eMkf����N�32p��)Q�M�;��5�q�fB��t&�gx�t���^s���������K�\vߺ1��i���N�AV��?h9&�p�1�3R{��#᧚]�ˏ��땪ALE OM0[�Xm�X%�����]��\`�P&eaP��~K#<_�e�KES;ԟ/�,���NF+W�VMQ�;�H�!������7'NZ�
۔J����`�hy-��݆��X�W�*]3H�)%��(Q��l�!ے�ŗ���K�,d��Jo��?TY�x��M�"���m״t��^��nl
���W�<ǌ|#D+b+��q2	��WaC\�li0-� �"�Bĉ�	����)��Х#�W�����q΂z�����]�`����zÂ�Yp��� !��H��o(�x��1�uU
P����(^�!�S}2��a������^W"�-��mv��N�/�)���kA���\��[g�$"\��>�0��5p�#��v+TZ�d�/n�0o����oe���-ֵb�Ee����j�VSқRx��H�/��]ٲi�:>]T�<}�2iHh�Zd܂���p�g��E�|]�����썵a�\�j`��-�A?�M0����N�_!J��!�4�Kz��:�Q��^�K��K(����]5q�`6��g�m���[�f�x���L-�%��ND|��*v�AMPج��R�v0���px����c,^�����t�6%s�C�ne���3y�'�,,�i����<.���������M u�jzp 9��\_a�Px�7����?�������ls<����u�XK�	S�Nu �\�n �3M�-�k3Ze���:��Gvj��\�A:U6Т]`hb��F�0�.����怹�q����6� �	\��R�b���|&0�kK=��0��X�J���d�����U��|j9��<�J�$��GFU~��xBx�+0G�����\�pO�4�z]��6����צ�H;�z�*�p��T�$�ĸ=�3�5ng��L�7�O��YlB}�������h�1�����`͆/h3x�����m.�}�d�����;��@#3�	���4F���l����p�y���HL�*C�Fh��=��4>�b����(�NU��E.e��λI=�d��x�8��!�$�X��v��QÀ�"���S{Ɏ��RT�q ��
��cޓ����/�$�q���K�Γ���V�UQt��~I\l�3_1)��C�	��U�܅!\+�Y�(��G�C��Z ͅ�"�r�/�
H�VZ�n�M�q? �5c�k��N[j��fț��xl�%�w8�~� �\ڱ3�2�̽��Í�VOA��-��O��)�����/���uJ��	)ɴ[;� ��"uk���l8F��>���9B���@糱%��(��Od�!��A���
OZ�l��H˪��z͠���$DL��E{�2���NG�?px�o�]z��Uf;NtM�b1u�N�KT�GNɠ��;x#uP��o?ߊ�Fy��"]����cR�-%E��6I�ߩ�S��:�+�S�JIn2��8BVU��gE����{�r���G{����#j�ȕ0��i�-6{H��E���':��4v��5��
g&m��`���� ���|���~� ���q:b�e�ϛ�׻}EK=�1��ʒ���v��������\�j�"��N�C(»�c�0[�`&ϡ���kF�Hv%��y>%<iFظ���N��t{��_T'*�d��8��������/㈙�F�/��)�B�f[�L�l3�U�UM�	O$}B���hv%B��&1��ӪUF�'�T�޷+�!���?���	D�k�-	S*�tOX^~:Fg�F�yl��'�Z�|�LCY�Fs�F�0o	\��~�i�%��հ
(!�.4��^T�W9�����B�`G�>��[�f}:;K�j��Xł�l�*l_�D�Hu����Cg�8�O���&�%��Y��s�_Lw�A���{�h��ƳT�p�I&� ���,��<�Cy���i3R�]{J.�T�Y[y�5��26g��Q7�@��E�?���'A��r���ű��F}y����	�+�N&��'�/K8�o�.�������G7��̬)^8���9�1<w0�NQoѨ)o�N�}��vy\ �J8"���<� �Kn��JnY\��f� �:H*K��y�1P�Ư;�u�6�(�����ڷ�}��p�SIП��4������;��x�"�|L�Fbq_f���`��I���_�30�d@4�ۦ#��&*���B�י���<�1\b6�kd�a��.ÐZpX��4�_�+>��<�1ß��H�uQ��[��ve[2�5�S�|��7$�V.�2lԹn�"��?)�R ����ѣ]Y1�z��W���<�yY,��f���y?ck+6��u��2/<�����?.D��2�x��(x0����R�&k��E_h��n�/�i9@�.e�[g�"�1��3,�
*P{DHċ2���S��4C�N� $��:&�*��\��O��@2bƟ�x蟌���q#ӊ�W�On�shGX������a�d�.V��&��s	�R�*�Eִ�Q���oDG%ޢ� "d��Ě���MX�����NI�1��.�ɍ-Dc࿁�XUth������sǝv&��Te�>��|n�,���p�@�vƗ�	\��������I8�� ^�N�G�r���Sx��C��Ͻ�!5�XAC�J�[-��&Z�ō+Ww��zE>�g��[����>����F�N��\.��N�w�:��9�YP:�L_v;��Y�C�O"siL9&���q�1܇T��򅙞+��|	L�E�g\�C:5o%8�*h�)�k��Lqh+P���0h�+OeIf�݊^b�����Ϫ�/ɓ��XV�Y9���RQ���:���@s#�)U�Ǳ-gI*�^��lH��f���ږt��bK�/��uʄ�AĶkf��<�,��*��$ ���S�RUT�>fͪy�����@�����-���^ &T����'�tO9pje ��?�J��5aђ�b�򨫭\*Vp8����N#�+xI��U���vo;y�I2$��)��#~�A`�洘vb7�gsq:�
2
ť:B����Arr"�|�VQ��e�a��DT�*EsNT�T�1�l<V���=7fꆷ�Zh#Ca�e2}_,�]��]�C�+����UĦ�|/jac_��4�G� 湓HV8��J�S
����켂�$�3���mHn�(g��P����.���s'Ϯ�K�Ѱ2�>�\����b)k;���%�-x��fzW�1�W&=���$�v?�7\e�H��rm�w\xZ��/o�B��C�]kD��eM�ӑƅ��"S�.2���	*��79�Fw��Ȝ��h�2B���i~ӷ�%W��x^�%��R%P�4�}��M�.C���Q&ɛ���[�$�-�t��1����>�w�!�IS�QTl(��.���f-d�x1�
�_��=��v��H��we'�&�()�cFf�Xf����iwD���Li*��G~��zD�5�����9�Շֲ4$�G�����'��X^,�=@U����r9Ff7U�٭O���r6Ҧ2W��Ǭ�3uͱst<Ru��\r�bH.ሎ��1��	�Ͳ��sQ�͍<ׂ���?�y,��z��t�wt�B�>�~���|`��-.pFd�^��5ܘ�p-���w��p�j؜.���񥉀�nLmB��)��8Lt{3�����~`�q�^ �%���������a�����E����w'ū~��[��d=��3� e�e��:I��#:Z'#�ż�nU�(N=��@;D��Q^
;
N^) %����B�+b`�~�sx˃G�R���Qd�S�y(��'y�LX���E~����'����:�Tz��rՈ^�t�)A+{m�
�̎�(����g`Ꜹ��C�/Y>�)�}��O�_��p:}Z>DTt���z4`��Eե&�*�T��-	w �H���ꩂmb��M[��U�G}W��2�I��hD��^��HY��}@��O�ף���T��P�2UstH�yfs6�9�8��7
G������_�ʕsC�h��G���崙3
�����ꍆ��y��#Z)�Ҟ�f�w��#}�h�P�4�W[��'ydZ$D�y��05�2$oM)��]�b�e����'�r� �`N<���B��S�yI7b7�ӎnjz�(�"�`}A�P�� ��o�}la��ɼ��ķN���xC)~�L?V�_- ���4�wV:�j�|Z/��}I��1�!H�N���N{�7S2&j�9��YH�h6���,�..T��~���hp�����e3�}_}1N�Q�b|̌��m+S�4aJf�x�tE��B�D�qr�K���0.�1�:�	�G^�x�Ko��l�n�&���3!N�qOI�[��3.YoN�"�r/�������v�9Ѓ���]z�YQ��)B���9U��3t�"p7q?7[	w`�zR��S��R`T���N� ��QpoX�)[�R��ژDF���ɧ��Đ��4��)o7�ħ}¬̽�{� �_%�[aS@r7�?"娹G��˭�^���΢} Q>�[i���r�y3�Y���!��a �dP���}k,����{�_����0�}$��so;Net�>������Q��$u&@���'��ںS���³��Y2pr��zP����G��X�uu�b�alr��q��xE�տ�FJ�,h�Y�c8�g���!W���iy��T�h�|a�xf9������tn��B����x3���ŭ�L�)�m���f�T����v@��E]v�9���vW�&�ڏ5yγ$^=R�jPQ)2<tP��2���٦��):�g$��Ӓ���(т��Ϋ��<G����/F���&����ݱ���>�X�*�k����h�F�g.g7�Ь1�ar�M�mξ���WpϦČb���|l��u\����fvQ{S�i�[�Mxcm�;G?��Ϝ��GF� �e�Q���Z�Ŭ�L�5�)��M&4�� G�բ�-� �1n�=�:jbW=1�h�"� �CG�ı۬u?��z���-GD�zM�S؎�TV�/]��T��וP���8��dOe�/�RwZQ^n��؁71�b�h��-i��2��j���E-��ƞ<�ÑfφL"v���{�1l�u�RABA�֔�u�5�:n�u�"�y|��hڋvlruj"S�3��x\MdÄ��*l���_W�A������B��f�P~�*���ȟ�_�J��K�σ�4��9l�3�tINtz�+�rma�c	x= ��r��6@�5m�K�����������sk�̟�'dc�V�M9�AZ�h�&�_��N��>(�s߆b :U+�W��C�$���4�C�o���F-!m�V�]��a�N2��l_��E�M��Y8�֍�1�Yg��n�8Q�YO�7,^�.�; ��Ӱ��-_Oy^��x�$�[a]xt��s}5�V8�#�&���5��3^���N{#W%�@ ��{�㺵j�l���?NnE�"�o�H?{�� �<%o�<l�{��E�f��������@�pg5e;A3��4&�wɌ���� ����&���j39�Q��Nd4@�0�7�'0}� �@w�ݠ��u�FHF$��5�I�ر��Z��J�K�k